module picorv32a (clk,
    mem_instr,
    mem_la_read,
    mem_la_write,
    mem_ready,
    mem_valid,
    pcpi_ready,
    pcpi_valid,
    pcpi_wait,
    pcpi_wr,
    resetn,
    trace_valid,
    trap,
    eoi,
    irq,
    mem_addr,
    mem_la_addr,
    mem_la_wdata,
    mem_la_wstrb,
    mem_rdata,
    mem_wdata,
    mem_wstrb,
    pcpi_insn,
    pcpi_rd,
    pcpi_rs1,
    pcpi_rs2,
    trace_data);
 input clk;
 output mem_instr;
 output mem_la_read;
 output mem_la_write;
 input mem_ready;
 output mem_valid;
 input pcpi_ready;
 output pcpi_valid;
 input pcpi_wait;
 input pcpi_wr;
 input resetn;
 output trace_valid;
 output trap;
 output [31:0] eoi;
 input [31:0] irq;
 output [31:0] mem_addr;
 output [31:0] mem_la_addr;
 output [31:0] mem_la_wdata;
 output [3:0] mem_la_wstrb;
 input [31:0] mem_rdata;
 output [31:0] mem_wdata;
 output [3:0] mem_wstrb;
 output [31:0] pcpi_insn;
 input [31:0] pcpi_rd;
 output [31:0] pcpi_rs1;
 output [31:0] pcpi_rs2;
 output [35:0] trace_data;

 sky130_vsdinv _20979_ (.A(net101),
    .Y(_18308_));
 sky130_fd_sc_hd__buf_4 _20980_ (.A(_18308_),
    .X(_18309_));
 sky130_fd_sc_hd__buf_4 _20981_ (.A(_18309_),
    .X(_18310_));
 sky130_fd_sc_hd__buf_2 _20982_ (.A(_18310_),
    .X(_18311_));
 sky130_fd_sc_hd__clkinv_4 _20983_ (.A(mem_do_prefetch),
    .Y(_18312_));
 sky130_fd_sc_hd__nand2_4 _20984_ (.A(net237),
    .B(net511),
    .Y(_18313_));
 sky130_vsdinv _20985_ (.A(_18313_),
    .Y(mem_xfer));
 sky130_vsdinv _20986_ (.A(\mem_state[1] ),
    .Y(_18314_));
 sky130_vsdinv _20987_ (.A(\mem_state[0] ),
    .Y(_18315_));
 sky130_fd_sc_hd__nor2_1 _20988_ (.A(_18314_),
    .B(_18315_),
    .Y(_18316_));
 sky130_fd_sc_hd__nor2_8 _20989_ (.A(\mem_state[1] ),
    .B(\mem_state[0] ),
    .Y(_00290_));
 sky130_vsdinv _20990_ (.A(_00290_),
    .Y(_18317_));
 sky130_fd_sc_hd__o21a_1 _20991_ (.A1(mem_xfer),
    .A2(_18316_),
    .B1(_18317_),
    .X(_18318_));
 sky130_fd_sc_hd__nor2_8 _20992_ (.A(mem_do_wdata),
    .B(mem_do_rdata),
    .Y(_18319_));
 sky130_vsdinv _20993_ (.A(mem_do_rinst),
    .Y(_18320_));
 sky130_fd_sc_hd__o21ai_2 _20994_ (.A1(_18313_),
    .A2(_18319_),
    .B1(_18320_),
    .Y(_18321_));
 sky130_fd_sc_hd__nand2_4 _20995_ (.A(_18318_),
    .B(_18321_),
    .Y(_18322_));
 sky130_vsdinv _20996_ (.A(_18322_),
    .Y(_18323_));
 sky130_fd_sc_hd__nor2_4 _20997_ (.A(_18312_),
    .B(_18323_),
    .Y(_18324_));
 sky130_fd_sc_hd__nor2_2 _20998_ (.A(_18311_),
    .B(_18324_),
    .Y(_18325_));
 sky130_vsdinv _20999_ (.A(mem_do_rdata),
    .Y(_18326_));
 sky130_vsdinv _21000_ (.A(\cpu_state[6] ),
    .Y(_18327_));
 sky130_fd_sc_hd__buf_2 _21001_ (.A(_18327_),
    .X(_18328_));
 sky130_fd_sc_hd__nor2_4 _21002_ (.A(_18326_),
    .B(_18328_),
    .Y(_00319_));
 sky130_fd_sc_hd__a21oi_4 _21003_ (.A1(_18325_),
    .A2(_00319_),
    .B1(_00332_),
    .Y(_18329_));
 sky130_fd_sc_hd__clkbuf_4 _21004_ (.A(net101),
    .X(_18330_));
 sky130_fd_sc_hd__buf_4 _21005_ (.A(_18330_),
    .X(_18331_));
 sky130_fd_sc_hd__buf_2 _21006_ (.A(_18331_),
    .X(_18332_));
 sky130_fd_sc_hd__clkbuf_4 _21007_ (.A(_18332_),
    .X(_18333_));
 sky130_fd_sc_hd__clkbuf_4 _21008_ (.A(\cpu_state[6] ),
    .X(_18334_));
 sky130_fd_sc_hd__a21bo_1 _21009_ (.A1(instr_lb),
    .A2(_18334_),
    .B1_N(_18329_),
    .X(_18335_));
 sky130_fd_sc_hd__o211a_1 _21010_ (.A1(latched_is_lb),
    .A2(_18329_),
    .B1(_18333_),
    .C1(_18335_),
    .X(_04071_));
 sky130_fd_sc_hd__clkbuf_4 _21011_ (.A(_18331_),
    .X(_18336_));
 sky130_fd_sc_hd__buf_4 _21012_ (.A(_18336_),
    .X(_18337_));
 sky130_fd_sc_hd__a21bo_1 _21013_ (.A1(instr_lh),
    .A2(_18334_),
    .B1_N(_18329_),
    .X(_18338_));
 sky130_fd_sc_hd__o211a_1 _21014_ (.A1(latched_is_lh),
    .A2(_18329_),
    .B1(_18337_),
    .C1(_18338_),
    .X(_04070_));
 sky130_vsdinv _21015_ (.A(instr_retirq),
    .Y(_18339_));
 sky130_fd_sc_hd__nand2_1 _21016_ (.A(_18339_),
    .B(net508),
    .Y(_18340_));
 sky130_vsdinv _21017_ (.A(_00331_),
    .Y(_18341_));
 sky130_fd_sc_hd__nand2_1 _21018_ (.A(_18340_),
    .B(_18341_),
    .Y(_18342_));
 sky130_vsdinv _21019_ (.A(latched_branch),
    .Y(_18343_));
 sky130_fd_sc_hd__clkbuf_4 _21020_ (.A(_18343_),
    .X(_18344_));
 sky130_fd_sc_hd__nand2_1 _21021_ (.A(_18342_),
    .B(_18344_),
    .Y(_18345_));
 sky130_fd_sc_hd__o211a_1 _21022_ (.A1(_20928_),
    .A2(_18342_),
    .B1(_18337_),
    .C1(_18345_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_4 _21023_ (.A(mem_do_rinst),
    .X(_18346_));
 sky130_fd_sc_hd__nor2_1 _21024_ (.A(_18346_),
    .B(mem_do_prefetch),
    .Y(_18347_));
 sky130_vsdinv _21025_ (.A(_18347_),
    .Y(_18348_));
 sky130_fd_sc_hd__nor2_1 _21026_ (.A(mem_do_rdata),
    .B(_18348_),
    .Y(_18349_));
 sky130_fd_sc_hd__inv_2 _21027_ (.A(mem_do_wdata),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_2 _21028_ (.A(_18349_),
    .B(_00291_),
    .Y(_18350_));
 sky130_fd_sc_hd__or2_1 _21029_ (.A(_18317_),
    .B(_18350_),
    .X(_18351_));
 sky130_vsdinv _21030_ (.A(net408),
    .Y(_18352_));
 sky130_fd_sc_hd__nor2_1 _21031_ (.A(\mem_state[0] ),
    .B(_18313_),
    .Y(_18353_));
 sky130_fd_sc_hd__a211o_1 _21032_ (.A1(\mem_state[0] ),
    .A2(_18346_),
    .B1(_18314_),
    .C1(_18353_),
    .X(_18354_));
 sky130_fd_sc_hd__a31o_1 _21033_ (.A1(_18351_),
    .A2(_18352_),
    .A3(_18354_),
    .B1(_18311_),
    .X(_18355_));
 sky130_fd_sc_hd__and2_1 _21034_ (.A(_18355_),
    .B(_00300_),
    .X(_18356_));
 sky130_fd_sc_hd__nor2_4 _21035_ (.A(net408),
    .B(_18310_),
    .Y(_18357_));
 sky130_fd_sc_hd__clkbuf_2 _21036_ (.A(_18357_),
    .X(_18358_));
 sky130_fd_sc_hd__nor2_1 _21037_ (.A(_18314_),
    .B(_18356_),
    .Y(_18359_));
 sky130_fd_sc_hd__a31o_1 _21038_ (.A1(_20893_),
    .A2(_18356_),
    .A3(_18358_),
    .B1(_18359_),
    .X(_04068_));
 sky130_fd_sc_hd__nor2_1 _21039_ (.A(_18315_),
    .B(_18356_),
    .Y(_18360_));
 sky130_fd_sc_hd__a31o_1 _21040_ (.A1(_20892_),
    .A2(_18356_),
    .A3(_18358_),
    .B1(_18360_),
    .X(_04067_));
 sky130_fd_sc_hd__nor2_4 _21041_ (.A(_18309_),
    .B(_18322_),
    .Y(_18361_));
 sky130_vsdinv _21042_ (.A(_18361_),
    .Y(_18362_));
 sky130_fd_sc_hd__nor2_1 _21043_ (.A(_18320_),
    .B(_18362_),
    .Y(_18363_));
 sky130_fd_sc_hd__buf_2 _21044_ (.A(_18363_),
    .X(_18364_));
 sky130_fd_sc_hd__clkbuf_4 _21045_ (.A(_18364_),
    .X(_20895_));
 sky130_fd_sc_hd__inv_2 _21046_ (.A(\decoded_rs1[4] ),
    .Y(_00366_));
 sky130_fd_sc_hd__clkbuf_2 _21047_ (.A(_18363_),
    .X(_18365_));
 sky130_fd_sc_hd__clkbuf_4 _21048_ (.A(_18365_),
    .X(_18366_));
 sky130_fd_sc_hd__or3_4 _21049_ (.A(\mem_rdata_latched[31] ),
    .B(\mem_rdata_latched[30] ),
    .C(\mem_rdata_latched[29] ),
    .X(_18367_));
 sky130_fd_sc_hd__or3_4 _21050_ (.A(\mem_rdata_latched[26] ),
    .B(\mem_rdata_latched[25] ),
    .C(_18367_),
    .X(_18368_));
 sky130_vsdinv _21051_ (.A(_00327_),
    .Y(_18369_));
 sky130_fd_sc_hd__or3_1 _21052_ (.A(\mem_rdata_latched[28] ),
    .B(_00330_),
    .C(_18369_),
    .X(_18370_));
 sky130_fd_sc_hd__and3b_1 _21053_ (.A_N(_00326_),
    .B(_00325_),
    .C(_00324_),
    .X(_18371_));
 sky130_fd_sc_hd__or4b_4 _21054_ (.A(_00329_),
    .B(_00328_),
    .C(_18370_),
    .D_N(_18371_),
    .X(_18372_));
 sky130_fd_sc_hd__nor2_1 _21055_ (.A(\mem_rdata_latched[27] ),
    .B(_18372_),
    .Y(_18373_));
 sky130_fd_sc_hd__and2b_1 _21056_ (.A_N(_18368_),
    .B(_18373_),
    .X(_18374_));
 sky130_fd_sc_hd__clkbuf_4 _21057_ (.A(_18364_),
    .X(_18375_));
 sky130_fd_sc_hd__o21ai_1 _21058_ (.A1(\mem_rdata_latched[19] ),
    .A2(_18374_),
    .B1(_18375_),
    .Y(_18376_));
 sky130_vsdinv _21059_ (.A(\mem_rdata_latched[25] ),
    .Y(_18377_));
 sky130_fd_sc_hd__and4b_1 _21060_ (.A_N(_18367_),
    .B(_18373_),
    .C(\mem_rdata_latched[26] ),
    .D(_18377_),
    .X(_18378_));
 sky130_fd_sc_hd__clkbuf_2 _21061_ (.A(_18378_),
    .X(_18379_));
 sky130_fd_sc_hd__nand2_1 _21062_ (.A(_18379_),
    .B(_18364_),
    .Y(_18380_));
 sky130_fd_sc_hd__o211ai_1 _21063_ (.A1(_00366_),
    .A2(_18366_),
    .B1(_18376_),
    .C1(_18380_),
    .Y(_04066_));
 sky130_fd_sc_hd__o21a_4 _21064_ (.A1(decoder_trigger),
    .A2(do_waitirq),
    .B1(instr_waitirq),
    .X(_00309_));
 sky130_vsdinv _21065_ (.A(decoder_trigger),
    .Y(_18381_));
 sky130_vsdinv _21066_ (.A(\irq_mask[6] ),
    .Y(_18382_));
 sky130_vsdinv _21067_ (.A(\irq_mask[4] ),
    .Y(_18383_));
 sky130_fd_sc_hd__and2_1 _21068_ (.A(_18383_),
    .B(\irq_pending[4] ),
    .X(_18384_));
 sky130_vsdinv _21069_ (.A(\irq_mask[5] ),
    .Y(_18385_));
 sky130_fd_sc_hd__and2_1 _21070_ (.A(_18385_),
    .B(\irq_pending[5] ),
    .X(_18386_));
 sky130_vsdinv _21071_ (.A(\irq_mask[7] ),
    .Y(_18387_));
 sky130_fd_sc_hd__and2_1 _21072_ (.A(_18387_),
    .B(\irq_pending[7] ),
    .X(_18388_));
 sky130_fd_sc_hd__a2111o_1 _21073_ (.A1(_18382_),
    .A2(\irq_pending[6] ),
    .B1(_18384_),
    .C1(_18386_),
    .D1(_18388_),
    .X(_18389_));
 sky130_vsdinv _21074_ (.A(\irq_mask[17] ),
    .Y(_18390_));
 sky130_fd_sc_hd__and2b_2 _21075_ (.A_N(\irq_mask[19] ),
    .B(\irq_pending[19] ),
    .X(_18391_));
 sky130_vsdinv _21076_ (.A(\irq_pending[16] ),
    .Y(_18392_));
 sky130_fd_sc_hd__nor2_4 _21077_ (.A(\irq_mask[16] ),
    .B(_18392_),
    .Y(_18393_));
 sky130_vsdinv _21078_ (.A(\irq_mask[18] ),
    .Y(_18394_));
 sky130_fd_sc_hd__and2_1 _21079_ (.A(_18394_),
    .B(\irq_pending[18] ),
    .X(_18395_));
 sky130_fd_sc_hd__a2111o_1 _21080_ (.A1(_18390_),
    .A2(\irq_pending[17] ),
    .B1(_18391_),
    .C1(_18393_),
    .D1(_18395_),
    .X(_18396_));
 sky130_vsdinv _21081_ (.A(\irq_mask[25] ),
    .Y(_18397_));
 sky130_vsdinv _21082_ (.A(\irq_mask[24] ),
    .Y(_18398_));
 sky130_fd_sc_hd__and2_1 _21083_ (.A(_18398_),
    .B(\irq_pending[24] ),
    .X(_18399_));
 sky130_vsdinv _21084_ (.A(\irq_mask[26] ),
    .Y(_18400_));
 sky130_fd_sc_hd__and2_1 _21085_ (.A(_18400_),
    .B(\irq_pending[26] ),
    .X(_18401_));
 sky130_vsdinv _21086_ (.A(\irq_mask[27] ),
    .Y(_18402_));
 sky130_fd_sc_hd__and2_1 _21087_ (.A(_18402_),
    .B(\irq_pending[27] ),
    .X(_18403_));
 sky130_fd_sc_hd__a2111o_1 _21088_ (.A1(_18397_),
    .A2(\irq_pending[25] ),
    .B1(_18399_),
    .C1(_18401_),
    .D1(_18403_),
    .X(_18404_));
 sky130_vsdinv _21089_ (.A(\irq_mask[10] ),
    .Y(_18405_));
 sky130_vsdinv _21090_ (.A(\irq_mask[8] ),
    .Y(_18406_));
 sky130_fd_sc_hd__and2b_1 _21091_ (.A_N(\irq_mask[9] ),
    .B(\irq_pending[9] ),
    .X(_18407_));
 sky130_vsdinv _21092_ (.A(\irq_mask[11] ),
    .Y(_18408_));
 sky130_fd_sc_hd__and2_1 _21093_ (.A(_18408_),
    .B(\irq_pending[11] ),
    .X(_18409_));
 sky130_fd_sc_hd__or2_1 _21094_ (.A(_18407_),
    .B(_18409_),
    .X(_18410_));
 sky130_fd_sc_hd__a221o_1 _21095_ (.A1(_18405_),
    .A2(\irq_pending[10] ),
    .B1(_18406_),
    .B2(\irq_pending[8] ),
    .C1(_18410_),
    .X(_18411_));
 sky130_fd_sc_hd__or4_4 _21096_ (.A(_18389_),
    .B(_18396_),
    .C(_18404_),
    .D(_18411_),
    .X(_18412_));
 sky130_vsdinv _21097_ (.A(\irq_mask[2] ),
    .Y(_18413_));
 sky130_vsdinv _21098_ (.A(\irq_pending[0] ),
    .Y(_18414_));
 sky130_fd_sc_hd__nor2_4 _21099_ (.A(\irq_mask[0] ),
    .B(_18414_),
    .Y(_18415_));
 sky130_vsdinv _21100_ (.A(\irq_pending[1] ),
    .Y(_18416_));
 sky130_fd_sc_hd__nor2_4 _21101_ (.A(\irq_mask[1] ),
    .B(_18416_),
    .Y(_18417_));
 sky130_vsdinv _21102_ (.A(\irq_mask[3] ),
    .Y(_18418_));
 sky130_fd_sc_hd__and2_1 _21103_ (.A(_18418_),
    .B(\irq_pending[3] ),
    .X(_18419_));
 sky130_fd_sc_hd__a2111o_1 _21104_ (.A1(_18413_),
    .A2(\irq_pending[2] ),
    .B1(_18415_),
    .C1(_18417_),
    .D1(_18419_),
    .X(_18420_));
 sky130_vsdinv _21105_ (.A(\irq_mask[21] ),
    .Y(_18421_));
 sky130_fd_sc_hd__and2b_2 _21106_ (.A_N(\irq_mask[22] ),
    .B(\irq_pending[22] ),
    .X(_18422_));
 sky130_vsdinv _21107_ (.A(\irq_mask[23] ),
    .Y(_18423_));
 sky130_fd_sc_hd__and2_1 _21108_ (.A(_18423_),
    .B(\irq_pending[23] ),
    .X(_18424_));
 sky130_vsdinv _21109_ (.A(\irq_mask[20] ),
    .Y(_18425_));
 sky130_fd_sc_hd__and2_1 _21110_ (.A(_18425_),
    .B(\irq_pending[20] ),
    .X(_18426_));
 sky130_fd_sc_hd__a2111o_2 _21111_ (.A1(_18421_),
    .A2(\irq_pending[21] ),
    .B1(_18422_),
    .C1(_18424_),
    .D1(_18426_),
    .X(_18427_));
 sky130_vsdinv _21112_ (.A(\irq_mask[14] ),
    .Y(_18428_));
 sky130_vsdinv _21113_ (.A(\irq_mask[12] ),
    .Y(_18429_));
 sky130_fd_sc_hd__and2b_2 _21114_ (.A_N(\irq_mask[13] ),
    .B(\irq_pending[13] ),
    .X(_18430_));
 sky130_fd_sc_hd__and2b_1 _21115_ (.A_N(\irq_mask[15] ),
    .B(\irq_pending[15] ),
    .X(_18431_));
 sky130_fd_sc_hd__or2_1 _21116_ (.A(_18430_),
    .B(_18431_),
    .X(_18432_));
 sky130_fd_sc_hd__a221o_1 _21117_ (.A1(_18428_),
    .A2(\irq_pending[14] ),
    .B1(_18429_),
    .B2(\irq_pending[12] ),
    .C1(_18432_),
    .X(_18433_));
 sky130_vsdinv _21118_ (.A(\irq_mask[30] ),
    .Y(_18434_));
 sky130_vsdinv _21119_ (.A(\irq_mask[28] ),
    .Y(_18435_));
 sky130_vsdinv _21120_ (.A(\irq_mask[29] ),
    .Y(_18436_));
 sky130_fd_sc_hd__and2_1 _21121_ (.A(_18436_),
    .B(\irq_pending[29] ),
    .X(_18437_));
 sky130_vsdinv _21122_ (.A(\irq_mask[31] ),
    .Y(_18438_));
 sky130_fd_sc_hd__and2_1 _21123_ (.A(_18438_),
    .B(\irq_pending[31] ),
    .X(_18439_));
 sky130_fd_sc_hd__or2_1 _21124_ (.A(_18437_),
    .B(_18439_),
    .X(_18440_));
 sky130_fd_sc_hd__a221o_1 _21125_ (.A1(_18434_),
    .A2(\irq_pending[30] ),
    .B1(_18435_),
    .B2(\irq_pending[28] ),
    .C1(_18440_),
    .X(_18441_));
 sky130_fd_sc_hd__or4_4 _21126_ (.A(_18420_),
    .B(_18427_),
    .C(_18433_),
    .D(_18441_),
    .X(_18442_));
 sky130_fd_sc_hd__nor2_1 _21127_ (.A(_18412_),
    .B(_18442_),
    .Y(_18443_));
 sky130_fd_sc_hd__or4_4 _21128_ (.A(irq_active),
    .B(irq_delay),
    .C(_18381_),
    .D(_18443_),
    .X(_18444_));
 sky130_fd_sc_hd__nor2_1 _21129_ (.A(\irq_state[1] ),
    .B(\irq_state[0] ),
    .Y(_18445_));
 sky130_fd_sc_hd__nand2_2 _21130_ (.A(_18444_),
    .B(_18445_),
    .Y(_18446_));
 sky130_fd_sc_hd__nor2_1 _21131_ (.A(_00309_),
    .B(_18446_),
    .Y(_18447_));
 sky130_fd_sc_hd__and3_4 _21132_ (.A(_18447_),
    .B(\cpu_state[1] ),
    .C(decoder_trigger),
    .X(_18448_));
 sky130_vsdinv _21133_ (.A(irq_active),
    .Y(_18449_));
 sky130_fd_sc_hd__nand2_1 _21134_ (.A(_18448_),
    .B(_18449_),
    .Y(_18450_));
 sky130_fd_sc_hd__o211a_1 _21135_ (.A1(irq_delay),
    .A2(_18448_),
    .B1(_18337_),
    .C1(_18450_),
    .X(_04065_));
 sky130_fd_sc_hd__buf_4 _21136_ (.A(net330),
    .X(_18451_));
 sky130_vsdinv _21137_ (.A(net291),
    .Y(_18452_));
 sky130_fd_sc_hd__or4_4 _21138_ (.A(net293),
    .B(net292),
    .C(net279),
    .D(_18452_),
    .X(_18453_));
 sky130_fd_sc_hd__nand2_2 _21139_ (.A(_18330_),
    .B(net370),
    .Y(_18454_));
 sky130_fd_sc_hd__or4_4 _21140_ (.A(net298),
    .B(net297),
    .C(net295),
    .D(net294),
    .X(_18455_));
 sky130_fd_sc_hd__nor2_2 _21141_ (.A(_18454_),
    .B(_18455_),
    .Y(_18456_));
 sky130_vsdinv _21142_ (.A(net302),
    .Y(_18457_));
 sky130_fd_sc_hd__and4b_1 _21143_ (.A_N(net299),
    .B(_18457_),
    .C(net301),
    .D(net300),
    .X(_18458_));
 sky130_fd_sc_hd__and3b_1 _21144_ (.A_N(net296),
    .B(net285),
    .C(net274),
    .X(_18459_));
 sky130_fd_sc_hd__and4b_1 _21145_ (.A_N(_18453_),
    .B(_18456_),
    .C(_18458_),
    .D(_18459_),
    .X(_18460_));
 sky130_vsdinv _21146_ (.A(\pcpi_mul.active[0] ),
    .Y(_18461_));
 sky130_vsdinv _21147_ (.A(\pcpi_mul.active[1] ),
    .Y(_18462_));
 sky130_fd_sc_hd__and3_4 _21148_ (.A(_18460_),
    .B(_18461_),
    .C(_18462_),
    .X(_18463_));
 sky130_fd_sc_hd__buf_4 _21149_ (.A(_18463_),
    .X(_18464_));
 sky130_fd_sc_hd__clkbuf_2 _21150_ (.A(_18464_),
    .X(_03728_));
 sky130_fd_sc_hd__or2_1 _21151_ (.A(net278),
    .B(net277),
    .X(_18465_));
 sky130_fd_sc_hd__nand2_1 _21152_ (.A(net278),
    .B(net277),
    .Y(_18466_));
 sky130_fd_sc_hd__buf_6 _21153_ (.A(\pcpi_mul.rs1[32] ),
    .X(_18467_));
 sky130_vsdinv _21154_ (.A(_18467_),
    .Y(_18468_));
 sky130_fd_sc_hd__buf_2 _21155_ (.A(_18468_),
    .X(_18469_));
 sky130_fd_sc_hd__nor2_1 _21156_ (.A(net465),
    .B(_18464_),
    .Y(_18470_));
 sky130_fd_sc_hd__a41o_1 _21157_ (.A1(_18451_),
    .A2(_03728_),
    .A3(_18465_),
    .A4(_18466_),
    .B1(_18470_),
    .X(_04064_));
 sky130_fd_sc_hd__buf_4 _21158_ (.A(net362),
    .X(_18471_));
 sky130_vsdinv _21159_ (.A(net278),
    .Y(_18472_));
 sky130_vsdinv _21160_ (.A(\pcpi_mul.rs2[32] ),
    .Y(_18473_));
 sky130_fd_sc_hd__buf_6 _21161_ (.A(_18473_),
    .X(_18474_));
 sky130_fd_sc_hd__buf_2 _21162_ (.A(_18474_),
    .X(_18475_));
 sky130_fd_sc_hd__clkbuf_4 _21163_ (.A(_18475_),
    .X(_18476_));
 sky130_fd_sc_hd__nor2_1 _21164_ (.A(_18476_),
    .B(_18464_),
    .Y(_18477_));
 sky130_fd_sc_hd__a41o_1 _21165_ (.A1(_18471_),
    .A2(_18472_),
    .A3(net277),
    .A4(_03728_),
    .B1(_18477_),
    .X(_04063_));
 sky130_fd_sc_hd__buf_2 _21166_ (.A(\cpu_state[4] ),
    .X(_18478_));
 sky130_fd_sc_hd__clkbuf_2 _21167_ (.A(_18478_),
    .X(_18479_));
 sky130_vsdinv _21168_ (.A(_00333_),
    .Y(_18480_));
 sky130_vsdinv _21169_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .Y(_18481_));
 sky130_fd_sc_hd__nor2_2 _21170_ (.A(alu_wait),
    .B(_18481_),
    .Y(_18482_));
 sky130_fd_sc_hd__nor2_1 _21171_ (.A(_18480_),
    .B(_18482_),
    .Y(_18483_));
 sky130_fd_sc_hd__clkbuf_4 _21172_ (.A(_18336_),
    .X(_18484_));
 sky130_fd_sc_hd__o221a_1 _21173_ (.A1(_18479_),
    .A2(_18480_),
    .B1(latched_stalu),
    .B2(_18483_),
    .C1(_18484_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_2 _21174_ (.A(latched_store),
    .X(_18485_));
 sky130_fd_sc_hd__buf_4 _21175_ (.A(_18485_),
    .X(_18486_));
 sky130_vsdinv _21176_ (.A(\cpu_state[4] ),
    .Y(_18487_));
 sky130_fd_sc_hd__inv_2 _21177_ (.A(alu_wait),
    .Y(_00302_));
 sky130_fd_sc_hd__or4_4 _21178_ (.A(instr_rdinstrh),
    .B(instr_rdinstr),
    .C(instr_rdcycleh),
    .D(instr_rdcycle),
    .X(_18488_));
 sky130_fd_sc_hd__nor2_2 _21179_ (.A(instr_setq),
    .B(instr_getq),
    .Y(_18489_));
 sky130_fd_sc_hd__nand2_2 _21180_ (.A(_18489_),
    .B(_18339_),
    .Y(_18490_));
 sky130_vsdinv _21181_ (.A(_18490_),
    .Y(_18491_));
 sky130_vsdinv _21182_ (.A(instr_timer),
    .Y(_18492_));
 sky130_fd_sc_hd__buf_2 _21183_ (.A(instr_maskirq),
    .X(_18493_));
 sky130_vsdinv _21184_ (.A(_18493_),
    .Y(_18494_));
 sky130_fd_sc_hd__and3_4 _21185_ (.A(_18491_),
    .B(_18492_),
    .C(_18494_),
    .X(_01717_));
 sky130_fd_sc_hd__and2b_1 _21186_ (.A_N(_18488_),
    .B(_01717_),
    .X(_18495_));
 sky130_fd_sc_hd__buf_4 _21187_ (.A(net508),
    .X(_18496_));
 sky130_fd_sc_hd__nand2_1 _21188_ (.A(_18495_),
    .B(_18496_),
    .Y(_18497_));
 sky130_fd_sc_hd__nor2_8 _21189_ (.A(net508),
    .B(\cpu_state[3] ),
    .Y(_18498_));
 sky130_fd_sc_hd__and3_1 _21190_ (.A(_18498_),
    .B(_18487_),
    .C(_18327_),
    .X(_18499_));
 sky130_fd_sc_hd__buf_4 _21191_ (.A(_18499_),
    .X(_01706_));
 sky130_vsdinv _21192_ (.A(\cpu_state[1] ),
    .Y(_18500_));
 sky130_fd_sc_hd__buf_2 _21193_ (.A(_18500_),
    .X(_18501_));
 sky130_fd_sc_hd__nand2_1 _21194_ (.A(_01706_),
    .B(_18501_),
    .Y(_18502_));
 sky130_fd_sc_hd__nor2_8 _21195_ (.A(instr_auipc),
    .B(instr_lui),
    .Y(_18503_));
 sky130_fd_sc_hd__inv_2 _21196_ (.A(instr_jal),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _21197_ (.A(_18503_),
    .B(_00323_),
    .Y(_00005_));
 sky130_fd_sc_hd__or4_4 _21198_ (.A(instr_sh),
    .B(instr_sb),
    .C(instr_lhu),
    .D(instr_lbu),
    .X(_18504_));
 sky130_fd_sc_hd__or4_1 _21199_ (.A(instr_lw),
    .B(instr_lh),
    .C(instr_lb),
    .D(instr_jalr),
    .X(_18505_));
 sky130_fd_sc_hd__or4_4 _21200_ (.A(instr_sra),
    .B(instr_srl),
    .C(instr_srai),
    .D(instr_srli),
    .X(_18506_));
 sky130_fd_sc_hd__or4_1 _21201_ (.A(_00005_),
    .B(_18504_),
    .C(_18505_),
    .D(_18506_),
    .X(_18507_));
 sky130_fd_sc_hd__or4_4 _21202_ (.A(instr_bltu),
    .B(instr_blt),
    .C(instr_bne),
    .D(instr_beq),
    .X(_18508_));
 sky130_fd_sc_hd__or4_4 _21203_ (.A(instr_andi),
    .B(instr_ori),
    .C(instr_xori),
    .D(instr_addi),
    .X(_18509_));
 sky130_fd_sc_hd__or4_4 _21204_ (.A(instr_slt),
    .B(instr_sll),
    .C(instr_sub),
    .D(instr_add),
    .X(_18510_));
 sky130_fd_sc_hd__or4_4 _21205_ (.A(instr_timer),
    .B(instr_waitirq),
    .C(instr_slli),
    .D(instr_sw),
    .X(_18511_));
 sky130_fd_sc_hd__or4_4 _21206_ (.A(_18508_),
    .B(_18509_),
    .C(_18510_),
    .D(_18511_),
    .X(_18512_));
 sky130_fd_sc_hd__or2_2 _21207_ (.A(_18507_),
    .B(_18512_),
    .X(_18513_));
 sky130_fd_sc_hd__or2_1 _21208_ (.A(instr_sltiu),
    .B(instr_slti),
    .X(_18514_));
 sky130_fd_sc_hd__or4_4 _21209_ (.A(instr_and),
    .B(instr_or),
    .C(instr_xor),
    .D(instr_sltu),
    .X(_18515_));
 sky130_fd_sc_hd__nor2_1 _21210_ (.A(instr_bgeu),
    .B(instr_bge),
    .Y(_18516_));
 sky130_fd_sc_hd__or3b_4 _21211_ (.A(_18514_),
    .B(_18515_),
    .C_N(_18516_),
    .X(_18517_));
 sky130_fd_sc_hd__or4_4 _21212_ (.A(instr_maskirq),
    .B(_18488_),
    .C(_18490_),
    .D(_18517_),
    .X(_18518_));
 sky130_fd_sc_hd__nor2_4 _21213_ (.A(_18513_),
    .B(_18518_),
    .Y(_00310_));
 sky130_fd_sc_hd__buf_2 _21214_ (.A(\cpu_state[3] ),
    .X(_18519_));
 sky130_fd_sc_hd__clkinv_4 _21215_ (.A(_18519_),
    .Y(_18520_));
 sky130_fd_sc_hd__a21o_1 _21216_ (.A1(_00310_),
    .A2(\pcpi_mul.active[1] ),
    .B1(_18520_),
    .X(_18521_));
 sky130_fd_sc_hd__o2111a_1 _21217_ (.A1(_18487_),
    .A2(_00302_),
    .B1(_18497_),
    .C1(_18502_),
    .D1(_18521_),
    .X(_18522_));
 sky130_fd_sc_hd__or2b_1 _21218_ (.A(_20929_),
    .B_N(_18522_),
    .X(_18523_));
 sky130_fd_sc_hd__o211a_1 _21219_ (.A1(_18486_),
    .A2(_18522_),
    .B1(_18337_),
    .C1(_18523_),
    .X(_04061_));
 sky130_fd_sc_hd__nor2_1 _21220_ (.A(\irq_state[1] ),
    .B(_18501_),
    .Y(_18524_));
 sky130_fd_sc_hd__clkbuf_4 _21221_ (.A(\irq_state[0] ),
    .X(_18525_));
 sky130_fd_sc_hd__buf_2 _21222_ (.A(_18525_),
    .X(_18526_));
 sky130_fd_sc_hd__nand2_1 _21223_ (.A(_18524_),
    .B(_18526_),
    .Y(_18527_));
 sky130_fd_sc_hd__clkbuf_4 _21224_ (.A(_18501_),
    .X(_18528_));
 sky130_fd_sc_hd__buf_1 _21225_ (.A(\irq_state[1] ),
    .X(_18529_));
 sky130_fd_sc_hd__clkbuf_4 _21226_ (.A(_18529_),
    .X(_18530_));
 sky130_fd_sc_hd__nand2_1 _21227_ (.A(_18528_),
    .B(_18530_),
    .Y(_18531_));
 sky130_fd_sc_hd__buf_2 _21228_ (.A(_18310_),
    .X(_18532_));
 sky130_fd_sc_hd__buf_2 _21229_ (.A(_18532_),
    .X(_18533_));
 sky130_fd_sc_hd__buf_4 _21230_ (.A(_18533_),
    .X(_18534_));
 sky130_fd_sc_hd__a21oi_1 _21231_ (.A1(_18527_),
    .A2(_18531_),
    .B1(_18534_),
    .Y(_04060_));
 sky130_fd_sc_hd__buf_2 _21232_ (.A(_18501_),
    .X(_18535_));
 sky130_vsdinv _21233_ (.A(_18445_),
    .Y(_18536_));
 sky130_fd_sc_hd__or3_2 _21234_ (.A(_18535_),
    .B(_18536_),
    .C(_18444_),
    .X(_18537_));
 sky130_fd_sc_hd__nand2_1 _21235_ (.A(_18528_),
    .B(_18526_),
    .Y(_18538_));
 sky130_fd_sc_hd__a21oi_1 _21236_ (.A1(_18537_),
    .A2(_18538_),
    .B1(_18534_),
    .Y(_04059_));
 sky130_fd_sc_hd__nor2_8 _21237_ (.A(\cpu_state[4] ),
    .B(_18496_),
    .Y(_18539_));
 sky130_fd_sc_hd__clkinv_4 _21238_ (.A(_18539_),
    .Y(_02542_));
 sky130_fd_sc_hd__nor2_1 _21239_ (.A(_18519_),
    .B(_02542_),
    .Y(_00354_));
 sky130_fd_sc_hd__nor2_2 _21240_ (.A(alu_wait),
    .B(_18487_),
    .Y(_18540_));
 sky130_vsdinv _21241_ (.A(net508),
    .Y(_18541_));
 sky130_fd_sc_hd__clkbuf_4 _21242_ (.A(_18541_),
    .X(_18542_));
 sky130_fd_sc_hd__buf_2 _21243_ (.A(_18542_),
    .X(_18543_));
 sky130_vsdinv _21244_ (.A(is_lb_lh_lw_lbu_lhu),
    .Y(_18544_));
 sky130_fd_sc_hd__nor2_1 _21245_ (.A(_18544_),
    .B(_00310_),
    .Y(_18545_));
 sky130_fd_sc_hd__nor2_1 _21246_ (.A(_18543_),
    .B(_18545_),
    .Y(_18546_));
 sky130_vsdinv _21247_ (.A(_00310_),
    .Y(_18547_));
 sky130_fd_sc_hd__a21oi_1 _21248_ (.A1(is_sb_sh_sw),
    .A2(_18547_),
    .B1(_18521_),
    .Y(_18548_));
 sky130_fd_sc_hd__a2111o_1 _21249_ (.A1(_18501_),
    .A2(_00354_),
    .B1(_18540_),
    .C1(_18546_),
    .D1(_18548_),
    .X(_18549_));
 sky130_fd_sc_hd__nor2_4 _21250_ (.A(_18309_),
    .B(_18323_),
    .Y(_18550_));
 sky130_fd_sc_hd__buf_4 _21251_ (.A(\cpu_state[1] ),
    .X(_18551_));
 sky130_fd_sc_hd__or4_4 _21252_ (.A(_18551_),
    .B(\cpu_state[0] ),
    .C(_18496_),
    .D(_18519_),
    .X(_18552_));
 sky130_fd_sc_hd__nor2_4 _21253_ (.A(\cpu_state[6] ),
    .B(\cpu_state[5] ),
    .Y(_00297_));
 sky130_vsdinv _21254_ (.A(_00297_),
    .Y(_18553_));
 sky130_vsdinv _21255_ (.A(_18482_),
    .Y(_18554_));
 sky130_fd_sc_hd__or4_4 _21256_ (.A(_18532_),
    .B(_00343_),
    .C(_18553_),
    .D(_18554_),
    .X(_18555_));
 sky130_fd_sc_hd__nor2_1 _21257_ (.A(_18552_),
    .B(_18555_),
    .Y(_18556_));
 sky130_vsdinv _21258_ (.A(_18550_),
    .Y(_18557_));
 sky130_fd_sc_hd__nor3_2 _21259_ (.A(_00356_),
    .B(_18557_),
    .C(_18549_),
    .Y(_18558_));
 sky130_fd_sc_hd__a311o_1 _21260_ (.A1(_18346_),
    .A2(_18549_),
    .A3(_18550_),
    .B1(_18556_),
    .C1(_18558_),
    .X(_04058_));
 sky130_fd_sc_hd__nor2_1 _21261_ (.A(instr_retirq),
    .B(instr_jalr),
    .Y(_18559_));
 sky130_fd_sc_hd__nand2_1 _21262_ (.A(_18448_),
    .B(_00323_),
    .Y(_18560_));
 sky130_fd_sc_hd__nand2_1 _21263_ (.A(_18560_),
    .B(_18312_),
    .Y(_18561_));
 sky130_fd_sc_hd__o211a_1 _21264_ (.A1(_18559_),
    .A2(_18560_),
    .B1(_18550_),
    .C1(_18561_),
    .X(_04057_));
 sky130_fd_sc_hd__nor2_1 _21265_ (.A(_00358_),
    .B(_00357_),
    .Y(_18562_));
 sky130_fd_sc_hd__nor2_1 _21266_ (.A(net493),
    .B(net491),
    .Y(_18563_));
 sky130_fd_sc_hd__and3_1 _21267_ (.A(_18562_),
    .B(_18563_),
    .C(_00368_),
    .X(_18564_));
 sky130_fd_sc_hd__buf_6 _21268_ (.A(_18564_),
    .X(_18565_));
 sky130_fd_sc_hd__nor2_8 _21269_ (.A(_01207_),
    .B(net437),
    .Y(\cpuregs_rs1[31] ));
 sky130_fd_sc_hd__nor2_4 _21270_ (.A(_18494_),
    .B(_18542_),
    .Y(_18566_));
 sky130_fd_sc_hd__clkbuf_2 _21271_ (.A(_18566_),
    .X(_18567_));
 sky130_fd_sc_hd__buf_2 _21272_ (.A(_18567_),
    .X(_18568_));
 sky130_fd_sc_hd__buf_4 _21273_ (.A(_18533_),
    .X(_18569_));
 sky130_fd_sc_hd__clkbuf_2 _21274_ (.A(_18567_),
    .X(_18570_));
 sky130_fd_sc_hd__nor2_1 _21275_ (.A(_18438_),
    .B(_18570_),
    .Y(_18571_));
 sky130_fd_sc_hd__a211o_1 _21276_ (.A1(\cpuregs_rs1[31] ),
    .A2(_18568_),
    .B1(_18569_),
    .C1(_18571_),
    .X(_04056_));
 sky130_vsdinv _21277_ (.A(_18566_),
    .Y(_18572_));
 sky130_fd_sc_hd__clkbuf_2 _21278_ (.A(_18572_),
    .X(_18573_));
 sky130_fd_sc_hd__buf_6 _21279_ (.A(_18564_),
    .X(_18574_));
 sky130_fd_sc_hd__nor2_2 _21280_ (.A(_18574_),
    .B(_18572_),
    .Y(_18575_));
 sky130_fd_sc_hd__clkbuf_2 _21281_ (.A(_18575_),
    .X(_18576_));
 sky130_vsdinv _21282_ (.A(_01180_),
    .Y(_18577_));
 sky130_fd_sc_hd__clkbuf_4 _21283_ (.A(_18310_),
    .X(_18578_));
 sky130_fd_sc_hd__buf_2 _21284_ (.A(_18578_),
    .X(_18579_));
 sky130_fd_sc_hd__a221o_1 _21285_ (.A1(\irq_mask[30] ),
    .A2(_18573_),
    .B1(_18576_),
    .B2(_18577_),
    .C1(_18579_),
    .X(_04055_));
 sky130_fd_sc_hd__buf_6 _21286_ (.A(_18574_),
    .X(_18580_));
 sky130_fd_sc_hd__nor2_8 _21287_ (.A(_01180_),
    .B(net427),
    .Y(\cpuregs_rs1[30] ));
 sky130_fd_sc_hd__buf_4 _21288_ (.A(_18574_),
    .X(_18581_));
 sky130_fd_sc_hd__nor2_8 _21289_ (.A(_01153_),
    .B(net426),
    .Y(\cpuregs_rs1[29] ));
 sky130_fd_sc_hd__nor2_1 _21290_ (.A(_18436_),
    .B(_18570_),
    .Y(_18582_));
 sky130_fd_sc_hd__a211o_1 _21291_ (.A1(\cpuregs_rs1[29] ),
    .A2(_18568_),
    .B1(_18569_),
    .C1(_18582_),
    .X(_04054_));
 sky130_vsdinv _21292_ (.A(_01126_),
    .Y(_18583_));
 sky130_fd_sc_hd__a221o_1 _21293_ (.A1(\irq_mask[28] ),
    .A2(_18573_),
    .B1(_18576_),
    .B2(_18583_),
    .C1(_18579_),
    .X(_04053_));
 sky130_fd_sc_hd__nor2_8 _21294_ (.A(_01126_),
    .B(net427),
    .Y(\cpuregs_rs1[28] ));
 sky130_vsdinv _21295_ (.A(_01099_),
    .Y(_18584_));
 sky130_fd_sc_hd__a221o_1 _21296_ (.A1(\irq_mask[27] ),
    .A2(_18573_),
    .B1(_18576_),
    .B2(_18584_),
    .C1(_18579_),
    .X(_04052_));
 sky130_fd_sc_hd__nor2_8 _21297_ (.A(_01099_),
    .B(net427),
    .Y(\cpuregs_rs1[27] ));
 sky130_fd_sc_hd__nor2_8 _21298_ (.A(_01072_),
    .B(net437),
    .Y(\cpuregs_rs1[26] ));
 sky130_fd_sc_hd__clkbuf_2 _21299_ (.A(_18567_),
    .X(_18585_));
 sky130_fd_sc_hd__nor2_1 _21300_ (.A(_18400_),
    .B(_18585_),
    .Y(_18586_));
 sky130_fd_sc_hd__a211o_1 _21301_ (.A1(\cpuregs_rs1[26] ),
    .A2(_18568_),
    .B1(_18569_),
    .C1(_18586_),
    .X(_04051_));
 sky130_fd_sc_hd__nor2_8 _21302_ (.A(_01045_),
    .B(net426),
    .Y(\cpuregs_rs1[25] ));
 sky130_fd_sc_hd__nor2_1 _21303_ (.A(_18397_),
    .B(_18585_),
    .Y(_18587_));
 sky130_fd_sc_hd__a211o_1 _21304_ (.A1(\cpuregs_rs1[25] ),
    .A2(_18568_),
    .B1(_18569_),
    .C1(_18587_),
    .X(_04050_));
 sky130_fd_sc_hd__nor2_8 _21305_ (.A(_01018_),
    .B(net437),
    .Y(\cpuregs_rs1[24] ));
 sky130_fd_sc_hd__nor2_1 _21306_ (.A(_18398_),
    .B(_18585_),
    .Y(_18588_));
 sky130_fd_sc_hd__a211o_1 _21307_ (.A1(\cpuregs_rs1[24] ),
    .A2(_18568_),
    .B1(_18569_),
    .C1(_18588_),
    .X(_04049_));
 sky130_fd_sc_hd__nor2_8 _21308_ (.A(_00991_),
    .B(net426),
    .Y(\cpuregs_rs1[23] ));
 sky130_fd_sc_hd__buf_4 _21309_ (.A(_18532_),
    .X(_18589_));
 sky130_fd_sc_hd__clkbuf_2 _21310_ (.A(_18589_),
    .X(_18590_));
 sky130_fd_sc_hd__nor2_1 _21311_ (.A(_18423_),
    .B(_18585_),
    .Y(_18591_));
 sky130_fd_sc_hd__a211o_1 _21312_ (.A1(\cpuregs_rs1[23] ),
    .A2(_18568_),
    .B1(_18590_),
    .C1(_18591_),
    .X(_04048_));
 sky130_vsdinv _21313_ (.A(_00964_),
    .Y(_18592_));
 sky130_fd_sc_hd__a221o_1 _21314_ (.A1(\irq_mask[22] ),
    .A2(_18573_),
    .B1(_18576_),
    .B2(_18592_),
    .C1(_18579_),
    .X(_04047_));
 sky130_fd_sc_hd__nor2_8 _21315_ (.A(_00964_),
    .B(net426),
    .Y(\cpuregs_rs1[22] ));
 sky130_vsdinv _21316_ (.A(_00937_),
    .Y(_18593_));
 sky130_fd_sc_hd__a221o_1 _21317_ (.A1(\irq_mask[21] ),
    .A2(_18573_),
    .B1(_18576_),
    .B2(_18593_),
    .C1(_18579_),
    .X(_04046_));
 sky130_fd_sc_hd__nor2_8 _21318_ (.A(_00937_),
    .B(_18580_),
    .Y(\cpuregs_rs1[21] ));
 sky130_fd_sc_hd__nor2_8 _21319_ (.A(_00910_),
    .B(net437),
    .Y(\cpuregs_rs1[20] ));
 sky130_fd_sc_hd__clkbuf_2 _21320_ (.A(_18567_),
    .X(_18594_));
 sky130_fd_sc_hd__nor2_1 _21321_ (.A(_18425_),
    .B(_18585_),
    .Y(_18595_));
 sky130_fd_sc_hd__a211o_1 _21322_ (.A1(\cpuregs_rs1[20] ),
    .A2(_18594_),
    .B1(_18590_),
    .C1(_18595_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_2 _21323_ (.A(_18572_),
    .X(_18596_));
 sky130_vsdinv _21324_ (.A(_00883_),
    .Y(_18597_));
 sky130_fd_sc_hd__buf_4 _21325_ (.A(_18578_),
    .X(_18598_));
 sky130_fd_sc_hd__a221o_1 _21326_ (.A1(\irq_mask[19] ),
    .A2(_18596_),
    .B1(_18576_),
    .B2(_18597_),
    .C1(_18598_),
    .X(_04044_));
 sky130_fd_sc_hd__nor2_8 _21327_ (.A(_00883_),
    .B(_18581_),
    .Y(\cpuregs_rs1[19] ));
 sky130_vsdinv _21328_ (.A(_00856_),
    .Y(_18599_));
 sky130_fd_sc_hd__a221o_1 _21329_ (.A1(\irq_mask[18] ),
    .A2(_18596_),
    .B1(_18575_),
    .B2(_18599_),
    .C1(_18598_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_8 _21330_ (.A(_00856_),
    .B(_18580_),
    .Y(\cpuregs_rs1[18] ));
 sky130_fd_sc_hd__buf_4 _21331_ (.A(_18574_),
    .X(_18600_));
 sky130_fd_sc_hd__nor2_8 _21332_ (.A(_00829_),
    .B(net425),
    .Y(\cpuregs_rs1[17] ));
 sky130_fd_sc_hd__nor2_1 _21333_ (.A(_18390_),
    .B(_18585_),
    .Y(_18601_));
 sky130_fd_sc_hd__a211o_1 _21334_ (.A1(\cpuregs_rs1[17] ),
    .A2(_18594_),
    .B1(_18590_),
    .C1(_18601_),
    .X(_04042_));
 sky130_vsdinv _21335_ (.A(_00802_),
    .Y(_18602_));
 sky130_fd_sc_hd__a221o_1 _21336_ (.A1(\irq_mask[16] ),
    .A2(_18596_),
    .B1(_18575_),
    .B2(_18602_),
    .C1(_18598_),
    .X(_04041_));
 sky130_fd_sc_hd__nor2_8 _21337_ (.A(_00802_),
    .B(_18581_),
    .Y(\cpuregs_rs1[16] ));
 sky130_fd_sc_hd__nor2_8 _21338_ (.A(_00775_),
    .B(_18565_),
    .Y(\cpuregs_rs1[15] ));
 sky130_vsdinv _21339_ (.A(\irq_mask[15] ),
    .Y(_18603_));
 sky130_fd_sc_hd__clkbuf_2 _21340_ (.A(_18567_),
    .X(_18604_));
 sky130_fd_sc_hd__nor2_1 _21341_ (.A(_18603_),
    .B(_18604_),
    .Y(_18605_));
 sky130_fd_sc_hd__a211o_1 _21342_ (.A1(\cpuregs_rs1[15] ),
    .A2(_18594_),
    .B1(_18590_),
    .C1(_18605_),
    .X(_04040_));
 sky130_fd_sc_hd__buf_4 _21343_ (.A(_18564_),
    .X(_18606_));
 sky130_fd_sc_hd__nor2_8 _21344_ (.A(_00748_),
    .B(net436),
    .Y(\cpuregs_rs1[14] ));
 sky130_fd_sc_hd__nor2_1 _21345_ (.A(_18428_),
    .B(_18604_),
    .Y(_18607_));
 sky130_fd_sc_hd__a211o_1 _21346_ (.A1(\cpuregs_rs1[14] ),
    .A2(_18594_),
    .B1(_18590_),
    .C1(_18607_),
    .X(_04039_));
 sky130_fd_sc_hd__nor2_8 _21347_ (.A(_00721_),
    .B(net425),
    .Y(\cpuregs_rs1[13] ));
 sky130_fd_sc_hd__and2_1 _21348_ (.A(_18596_),
    .B(\irq_mask[13] ),
    .X(_18608_));
 sky130_fd_sc_hd__a211o_1 _21349_ (.A1(\cpuregs_rs1[13] ),
    .A2(_18594_),
    .B1(_18590_),
    .C1(_18608_),
    .X(_04038_));
 sky130_fd_sc_hd__nor2_8 _21350_ (.A(_00694_),
    .B(net425),
    .Y(\cpuregs_rs1[12] ));
 sky130_fd_sc_hd__buf_2 _21351_ (.A(_18589_),
    .X(_18609_));
 sky130_fd_sc_hd__nor2_1 _21352_ (.A(_18429_),
    .B(_18604_),
    .Y(_18610_));
 sky130_fd_sc_hd__a211o_1 _21353_ (.A1(\cpuregs_rs1[12] ),
    .A2(_18594_),
    .B1(_18609_),
    .C1(_18610_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_8 _21354_ (.A(_00667_),
    .B(net436),
    .Y(\cpuregs_rs1[11] ));
 sky130_fd_sc_hd__clkbuf_2 _21355_ (.A(_18567_),
    .X(_18611_));
 sky130_fd_sc_hd__nor2_1 _21356_ (.A(_18408_),
    .B(_18604_),
    .Y(_18612_));
 sky130_fd_sc_hd__a211o_1 _21357_ (.A1(\cpuregs_rs1[11] ),
    .A2(_18611_),
    .B1(_18609_),
    .C1(_18612_),
    .X(_04036_));
 sky130_fd_sc_hd__nor2_8 _21358_ (.A(_00640_),
    .B(net436),
    .Y(\cpuregs_rs1[10] ));
 sky130_fd_sc_hd__nor2_1 _21359_ (.A(_18405_),
    .B(_18604_),
    .Y(_18613_));
 sky130_fd_sc_hd__a211o_1 _21360_ (.A1(\cpuregs_rs1[10] ),
    .A2(_18611_),
    .B1(_18609_),
    .C1(_18613_),
    .X(_04035_));
 sky130_fd_sc_hd__nor2_8 _21361_ (.A(_00613_),
    .B(net425),
    .Y(\cpuregs_rs1[9] ));
 sky130_fd_sc_hd__and2_1 _21362_ (.A(_18572_),
    .B(\irq_mask[9] ),
    .X(_18614_));
 sky130_fd_sc_hd__a211o_1 _21363_ (.A1(\cpuregs_rs1[9] ),
    .A2(_18611_),
    .B1(_18609_),
    .C1(_18614_),
    .X(_04034_));
 sky130_fd_sc_hd__nor2_8 _21364_ (.A(_00586_),
    .B(net436),
    .Y(\cpuregs_rs1[8] ));
 sky130_fd_sc_hd__nor2_1 _21365_ (.A(_18406_),
    .B(_18604_),
    .Y(_18615_));
 sky130_fd_sc_hd__a211o_1 _21366_ (.A1(\cpuregs_rs1[8] ),
    .A2(_18611_),
    .B1(_18609_),
    .C1(_18615_),
    .X(_04033_));
 sky130_fd_sc_hd__nor2_8 _21367_ (.A(_00559_),
    .B(_18600_),
    .Y(\cpuregs_rs1[7] ));
 sky130_fd_sc_hd__clkbuf_2 _21368_ (.A(_18566_),
    .X(_18616_));
 sky130_fd_sc_hd__nor2_1 _21369_ (.A(_18387_),
    .B(_18616_),
    .Y(_18617_));
 sky130_fd_sc_hd__a211o_1 _21370_ (.A1(\cpuregs_rs1[7] ),
    .A2(_18611_),
    .B1(_18609_),
    .C1(_18617_),
    .X(_04032_));
 sky130_vsdinv _21371_ (.A(_00532_),
    .Y(_18618_));
 sky130_fd_sc_hd__a221o_1 _21372_ (.A1(\irq_mask[6] ),
    .A2(_18596_),
    .B1(_18575_),
    .B2(_18618_),
    .C1(_18598_),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_8 _21373_ (.A(_00532_),
    .B(_18565_),
    .Y(\cpuregs_rs1[6] ));
 sky130_fd_sc_hd__nor2_8 _21374_ (.A(_00505_),
    .B(_18600_),
    .Y(\cpuregs_rs1[5] ));
 sky130_fd_sc_hd__buf_2 _21375_ (.A(_18578_),
    .X(_18619_));
 sky130_fd_sc_hd__nor2_1 _21376_ (.A(_18385_),
    .B(_18616_),
    .Y(_18620_));
 sky130_fd_sc_hd__a211o_1 _21377_ (.A1(\cpuregs_rs1[5] ),
    .A2(_18611_),
    .B1(_18619_),
    .C1(_18620_),
    .X(_04030_));
 sky130_fd_sc_hd__nor2_8 _21378_ (.A(_00478_),
    .B(_18580_),
    .Y(\cpuregs_rs1[4] ));
 sky130_fd_sc_hd__nor2_1 _21379_ (.A(_18383_),
    .B(_18616_),
    .Y(_18621_));
 sky130_fd_sc_hd__a211o_1 _21380_ (.A1(\cpuregs_rs1[4] ),
    .A2(_18570_),
    .B1(_18619_),
    .C1(_18621_),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_8 _21381_ (.A(_00451_),
    .B(_18606_),
    .Y(\cpuregs_rs1[3] ));
 sky130_fd_sc_hd__nor2_1 _21382_ (.A(_18418_),
    .B(_18616_),
    .Y(_18622_));
 sky130_fd_sc_hd__a211o_1 _21383_ (.A1(\cpuregs_rs1[3] ),
    .A2(_18570_),
    .B1(_18619_),
    .C1(_18622_),
    .X(_04028_));
 sky130_fd_sc_hd__nor2_8 _21384_ (.A(_00424_),
    .B(_18606_),
    .Y(\cpuregs_rs1[2] ));
 sky130_fd_sc_hd__buf_2 _21385_ (.A(_18413_),
    .X(_18623_));
 sky130_fd_sc_hd__nor2_1 _21386_ (.A(_18623_),
    .B(_18616_),
    .Y(_18624_));
 sky130_fd_sc_hd__a211o_1 _21387_ (.A1(\cpuregs_rs1[2] ),
    .A2(_18570_),
    .B1(_18619_),
    .C1(_18624_),
    .X(_04027_));
 sky130_fd_sc_hd__nor2_8 _21388_ (.A(_00397_),
    .B(_18574_),
    .Y(\cpuregs_rs1[1] ));
 sky130_vsdinv _21389_ (.A(\irq_mask[1] ),
    .Y(_18625_));
 sky130_fd_sc_hd__nor2_1 _21390_ (.A(_18625_),
    .B(_18616_),
    .Y(_18626_));
 sky130_fd_sc_hd__a211o_1 _21391_ (.A1(\cpuregs_rs1[1] ),
    .A2(_18570_),
    .B1(_18619_),
    .C1(_18626_),
    .X(_04026_));
 sky130_vsdinv _21392_ (.A(_18574_),
    .Y(_18627_));
 sky130_fd_sc_hd__nand2_2 _21393_ (.A(_18627_),
    .B(_00370_),
    .Y(_18628_));
 sky130_fd_sc_hd__nor2_1 _21394_ (.A(_18596_),
    .B(_18628_),
    .Y(_18629_));
 sky130_fd_sc_hd__a211o_1 _21395_ (.A1(\irq_mask[0] ),
    .A2(_18573_),
    .B1(_18619_),
    .C1(_18629_),
    .X(_04025_));
 sky130_vsdinv _21396_ (.A(_18628_),
    .Y(\cpuregs_rs1[0] ));
 sky130_fd_sc_hd__clkbuf_2 _21397_ (.A(mem_do_wdata),
    .X(_18630_));
 sky130_fd_sc_hd__clkbuf_4 _21398_ (.A(_18347_),
    .X(_00301_));
 sky130_fd_sc_hd__nor2_1 _21399_ (.A(_18630_),
    .B(_00301_),
    .Y(_18631_));
 sky130_vsdinv _21400_ (.A(_18357_),
    .Y(_18632_));
 sky130_fd_sc_hd__nand2_2 _21401_ (.A(_18350_),
    .B(_00290_),
    .Y(_18633_));
 sky130_fd_sc_hd__nor2_8 _21402_ (.A(_18632_),
    .B(_18633_),
    .Y(_18634_));
 sky130_fd_sc_hd__buf_6 _21403_ (.A(_18634_),
    .X(_18635_));
 sky130_fd_sc_hd__mux2_1 _21404_ (.A0(net166),
    .A1(_18631_),
    .S(_18635_),
    .X(_04024_));
 sky130_vsdinv _21405_ (.A(_00328_),
    .Y(_18636_));
 sky130_fd_sc_hd__and3_1 _21406_ (.A(_18636_),
    .B(_00329_),
    .C(_00330_),
    .X(_18637_));
 sky130_vsdinv _21407_ (.A(_18365_),
    .Y(_18638_));
 sky130_fd_sc_hd__a31o_1 _21408_ (.A1(_18369_),
    .A2(_18371_),
    .A3(_18637_),
    .B1(_18638_),
    .X(_18639_));
 sky130_fd_sc_hd__o211a_1 _21409_ (.A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(_18366_),
    .B1(_18337_),
    .C1(_18639_),
    .X(_04023_));
 sky130_fd_sc_hd__nand2_2 _21410_ (.A(_18366_),
    .B(\mem_rdata_latched[18] ),
    .Y(_18640_));
 sky130_fd_sc_hd__clkbuf_4 _21411_ (.A(_18638_),
    .X(_00337_));
 sky130_fd_sc_hd__a2bb2o_1 _21412_ (.A1_N(_18640_),
    .A2_N(_18379_),
    .B1(\decoded_rs1[3] ),
    .B2(_00337_),
    .X(_04022_));
 sky130_fd_sc_hd__nand2_2 _21413_ (.A(_18375_),
    .B(\mem_rdata_latched[17] ),
    .Y(_18641_));
 sky130_fd_sc_hd__a2bb2o_1 _21414_ (.A1_N(_18641_),
    .A2_N(_18379_),
    .B1(\decoded_rs1[2] ),
    .B2(_00337_),
    .X(_04021_));
 sky130_fd_sc_hd__nand2_2 _21415_ (.A(_18375_),
    .B(\mem_rdata_latched[16] ),
    .Y(_18642_));
 sky130_fd_sc_hd__a2bb2o_1 _21416_ (.A1_N(_18642_),
    .A2_N(_18379_),
    .B1(\decoded_rs1[1] ),
    .B2(_00337_),
    .X(_04020_));
 sky130_fd_sc_hd__nand2_2 _21417_ (.A(_18375_),
    .B(\mem_rdata_latched[15] ),
    .Y(_18643_));
 sky130_fd_sc_hd__a2bb2o_1 _21418_ (.A1_N(_18643_),
    .A2_N(_18379_),
    .B1(\decoded_rs1[0] ),
    .B2(_00337_),
    .X(_04019_));
 sky130_fd_sc_hd__clkbuf_2 _21419_ (.A(_18533_),
    .X(_18644_));
 sky130_fd_sc_hd__nor2_2 _21420_ (.A(decoder_pseudo_trigger),
    .B(_18381_),
    .Y(_18645_));
 sky130_vsdinv _21421_ (.A(_18645_),
    .Y(_18646_));
 sky130_fd_sc_hd__clkbuf_4 _21422_ (.A(_18646_),
    .X(_18647_));
 sky130_fd_sc_hd__clkbuf_4 _21423_ (.A(_18647_),
    .X(_18648_));
 sky130_fd_sc_hd__inv_2 _21424_ (.A(\mem_rdata_q[14] ),
    .Y(_00334_));
 sky130_vsdinv _21425_ (.A(\mem_rdata_q[13] ),
    .Y(_18649_));
 sky130_fd_sc_hd__clkbuf_2 _21426_ (.A(_18649_),
    .X(_18650_));
 sky130_vsdinv _21427_ (.A(\mem_rdata_q[12] ),
    .Y(_18651_));
 sky130_fd_sc_hd__or3_4 _21428_ (.A(_00334_),
    .B(_18650_),
    .C(_18651_),
    .X(_18652_));
 sky130_vsdinv _21429_ (.A(is_alu_reg_reg),
    .Y(_18653_));
 sky130_fd_sc_hd__nor2_1 _21430_ (.A(\mem_rdata_q[28] ),
    .B(\mem_rdata_q[26] ),
    .Y(_18654_));
 sky130_vsdinv _21431_ (.A(\mem_rdata_q[27] ),
    .Y(_18655_));
 sky130_vsdinv _21432_ (.A(\mem_rdata_q[25] ),
    .Y(_18656_));
 sky130_fd_sc_hd__and3_1 _21433_ (.A(_18654_),
    .B(_18655_),
    .C(_18656_),
    .X(_18657_));
 sky130_vsdinv _21434_ (.A(\mem_rdata_q[31] ),
    .Y(_18658_));
 sky130_vsdinv _21435_ (.A(\mem_rdata_q[30] ),
    .Y(_18659_));
 sky130_vsdinv _21436_ (.A(\mem_rdata_q[29] ),
    .Y(_18660_));
 sky130_fd_sc_hd__and3_1 _21437_ (.A(_18658_),
    .B(_18659_),
    .C(_18660_),
    .X(_18661_));
 sky130_fd_sc_hd__and3_1 _21438_ (.A(_18657_),
    .B(_18661_),
    .C(_18645_),
    .X(_18662_));
 sky130_vsdinv _21439_ (.A(_18662_),
    .Y(_18663_));
 sky130_fd_sc_hd__nor2_4 _21440_ (.A(_18653_),
    .B(_18663_),
    .Y(_18664_));
 sky130_vsdinv _21441_ (.A(_18664_),
    .Y(_18665_));
 sky130_fd_sc_hd__o2bb2a_1 _21442_ (.A1_N(instr_and),
    .A2_N(_18648_),
    .B1(_18652_),
    .B2(_18665_),
    .X(_18666_));
 sky130_fd_sc_hd__nor2_1 _21443_ (.A(_18644_),
    .B(_18666_),
    .Y(_04018_));
 sky130_fd_sc_hd__buf_4 _21444_ (.A(\mem_rdata_q[14] ),
    .X(_18667_));
 sky130_fd_sc_hd__and3_1 _21445_ (.A(_18651_),
    .B(_18667_),
    .C(\mem_rdata_q[13] ),
    .X(_18668_));
 sky130_fd_sc_hd__nand2_1 _21446_ (.A(_18664_),
    .B(_18668_),
    .Y(_18669_));
 sky130_fd_sc_hd__clkbuf_4 _21447_ (.A(_18647_),
    .X(_18670_));
 sky130_fd_sc_hd__nand2_1 _21448_ (.A(_18670_),
    .B(instr_or),
    .Y(_18671_));
 sky130_fd_sc_hd__a21oi_1 _21449_ (.A1(_18669_),
    .A2(_18671_),
    .B1(_18534_),
    .Y(_04017_));
 sky130_fd_sc_hd__buf_2 _21450_ (.A(\mem_rdata_q[31] ),
    .X(_18672_));
 sky130_vsdinv _21451_ (.A(_18657_),
    .Y(_18673_));
 sky130_fd_sc_hd__nor2_1 _21452_ (.A(\mem_rdata_q[29] ),
    .B(_18646_),
    .Y(_18674_));
 sky130_vsdinv _21453_ (.A(_18674_),
    .Y(_18675_));
 sky130_fd_sc_hd__or4_4 _21454_ (.A(_18672_),
    .B(_18659_),
    .C(_18673_),
    .D(_18675_),
    .X(_18676_));
 sky130_vsdinv _21455_ (.A(_18676_),
    .Y(_18677_));
 sky130_fd_sc_hd__and3_1 _21456_ (.A(_18650_),
    .B(\mem_rdata_q[14] ),
    .C(\mem_rdata_q[12] ),
    .X(_18678_));
 sky130_vsdinv _21457_ (.A(_18678_),
    .Y(_18679_));
 sky130_fd_sc_hd__nor2_1 _21458_ (.A(_18653_),
    .B(_18679_),
    .Y(_18680_));
 sky130_fd_sc_hd__nand2_1 _21459_ (.A(_18677_),
    .B(_18680_),
    .Y(_18681_));
 sky130_fd_sc_hd__nand2_1 _21460_ (.A(_18670_),
    .B(instr_sra),
    .Y(_18682_));
 sky130_fd_sc_hd__buf_2 _21461_ (.A(_18533_),
    .X(_18683_));
 sky130_fd_sc_hd__a21oi_1 _21462_ (.A1(_18681_),
    .A2(_18682_),
    .B1(_18683_),
    .Y(_04016_));
 sky130_fd_sc_hd__buf_2 _21463_ (.A(_18662_),
    .X(_18684_));
 sky130_fd_sc_hd__nand2_1 _21464_ (.A(_18684_),
    .B(_18680_),
    .Y(_18685_));
 sky130_fd_sc_hd__nand2_1 _21465_ (.A(_18670_),
    .B(instr_srl),
    .Y(_18686_));
 sky130_fd_sc_hd__a21oi_1 _21466_ (.A1(_18685_),
    .A2(_18686_),
    .B1(_18683_),
    .Y(_04015_));
 sky130_fd_sc_hd__clkbuf_2 _21467_ (.A(_18646_),
    .X(_18687_));
 sky130_fd_sc_hd__and3_2 _21468_ (.A(_18650_),
    .B(_18651_),
    .C(_18667_),
    .X(_18688_));
 sky130_fd_sc_hd__a22o_1 _21469_ (.A1(instr_xor),
    .A2(_18687_),
    .B1(_18664_),
    .B2(_18688_),
    .X(_18689_));
 sky130_fd_sc_hd__and2_1 _21470_ (.A(_18689_),
    .B(_18484_),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_4 _21471_ (.A(_18646_),
    .X(_18690_));
 sky130_fd_sc_hd__and2_1 _21472_ (.A(_18690_),
    .B(instr_sltu),
    .X(_18691_));
 sky130_fd_sc_hd__clkbuf_4 _21473_ (.A(\mem_rdata_q[12] ),
    .X(_18692_));
 sky130_fd_sc_hd__nor2_2 _21474_ (.A(\mem_rdata_q[14] ),
    .B(_18650_),
    .Y(_18693_));
 sky130_fd_sc_hd__and3_1 _21475_ (.A(_18664_),
    .B(_18692_),
    .C(_18693_),
    .X(_18694_));
 sky130_fd_sc_hd__clkbuf_4 _21476_ (.A(_18331_),
    .X(_18695_));
 sky130_fd_sc_hd__clkbuf_4 _21477_ (.A(_18695_),
    .X(_18696_));
 sky130_fd_sc_hd__o21a_1 _21478_ (.A1(_18691_),
    .A2(_18694_),
    .B1(_18696_),
    .X(_04013_));
 sky130_fd_sc_hd__nand2_1 _21479_ (.A(_18693_),
    .B(_18651_),
    .Y(_18697_));
 sky130_vsdinv _21480_ (.A(_18697_),
    .Y(_18698_));
 sky130_fd_sc_hd__a22o_1 _21481_ (.A1(instr_slt),
    .A2(_18687_),
    .B1(_18664_),
    .B2(_18698_),
    .X(_18699_));
 sky130_fd_sc_hd__and2_1 _21482_ (.A(_18699_),
    .B(_18484_),
    .X(_04012_));
 sky130_fd_sc_hd__and3_2 _21483_ (.A(_00334_),
    .B(_18650_),
    .C(\mem_rdata_q[12] ),
    .X(_18700_));
 sky130_fd_sc_hd__a22o_1 _21484_ (.A1(instr_sll),
    .A2(_18687_),
    .B1(_18664_),
    .B2(_18700_),
    .X(_18701_));
 sky130_fd_sc_hd__and2_1 _21485_ (.A(_18701_),
    .B(_18484_),
    .X(_04011_));
 sky130_fd_sc_hd__and3_2 _21486_ (.A(_00334_),
    .B(_18649_),
    .C(_18651_),
    .X(_18702_));
 sky130_vsdinv _21487_ (.A(_18702_),
    .Y(_18703_));
 sky130_fd_sc_hd__or3_2 _21488_ (.A(_18653_),
    .B(_18703_),
    .C(_18676_),
    .X(_18704_));
 sky130_fd_sc_hd__nand2_1 _21489_ (.A(_18670_),
    .B(instr_sub),
    .Y(_18705_));
 sky130_fd_sc_hd__a21oi_1 _21490_ (.A1(_18704_),
    .A2(_18705_),
    .B1(_18683_),
    .Y(_04010_));
 sky130_fd_sc_hd__a32o_1 _21491_ (.A1(_18684_),
    .A2(is_alu_reg_reg),
    .A3(_18702_),
    .B1(instr_add),
    .B2(_18690_),
    .X(_18706_));
 sky130_fd_sc_hd__and2_1 _21492_ (.A(_18706_),
    .B(_18484_),
    .X(_04009_));
 sky130_vsdinv _21493_ (.A(decoder_pseudo_trigger),
    .Y(_18707_));
 sky130_fd_sc_hd__and3_2 _21494_ (.A(_18707_),
    .B(is_alu_reg_imm),
    .C(decoder_trigger),
    .X(_18708_));
 sky130_vsdinv _21495_ (.A(_18708_),
    .Y(_18709_));
 sky130_fd_sc_hd__o2bb2a_1 _21496_ (.A1_N(instr_andi),
    .A2_N(_18648_),
    .B1(_18709_),
    .B2(_18652_),
    .X(_18710_));
 sky130_fd_sc_hd__nor2_1 _21497_ (.A(_18644_),
    .B(_18710_),
    .Y(_04008_));
 sky130_fd_sc_hd__buf_2 _21498_ (.A(_18646_),
    .X(_18711_));
 sky130_fd_sc_hd__buf_2 _21499_ (.A(_18711_),
    .X(_18712_));
 sky130_fd_sc_hd__nand2_1 _21500_ (.A(_18712_),
    .B(instr_ori),
    .Y(_18713_));
 sky130_fd_sc_hd__nand2_1 _21501_ (.A(_18668_),
    .B(_18708_),
    .Y(_18714_));
 sky130_fd_sc_hd__a21oi_1 _21502_ (.A1(_18713_),
    .A2(_18714_),
    .B1(_18683_),
    .Y(_04007_));
 sky130_fd_sc_hd__a22o_1 _21503_ (.A1(_18688_),
    .A2(_18708_),
    .B1(_18690_),
    .B2(instr_xori),
    .X(_18715_));
 sky130_fd_sc_hd__and2_1 _21504_ (.A(_18715_),
    .B(_18484_),
    .X(_04006_));
 sky130_fd_sc_hd__and3_1 _21505_ (.A(_18708_),
    .B(_18692_),
    .C(_18693_),
    .X(_18716_));
 sky130_fd_sc_hd__and2_1 _21506_ (.A(_18687_),
    .B(instr_sltiu),
    .X(_18717_));
 sky130_fd_sc_hd__o21a_1 _21507_ (.A1(_18716_),
    .A2(_18717_),
    .B1(_18696_),
    .X(_04005_));
 sky130_fd_sc_hd__o2bb2a_1 _21508_ (.A1_N(instr_slti),
    .A2_N(_18648_),
    .B1(_18697_),
    .B2(_18709_),
    .X(_18718_));
 sky130_fd_sc_hd__nor2_1 _21509_ (.A(_18644_),
    .B(_18718_),
    .Y(_04004_));
 sky130_fd_sc_hd__a22o_1 _21510_ (.A1(_18702_),
    .A2(_18708_),
    .B1(instr_addi),
    .B2(_18690_),
    .X(_18719_));
 sky130_fd_sc_hd__and2_1 _21511_ (.A(_18719_),
    .B(_18333_),
    .X(_04003_));
 sky130_fd_sc_hd__nor2_4 _21512_ (.A(_18481_),
    .B(_18646_),
    .Y(_18720_));
 sky130_vsdinv _21513_ (.A(_18720_),
    .Y(_18721_));
 sky130_fd_sc_hd__o2bb2a_1 _21514_ (.A1_N(instr_bgeu),
    .A2_N(_18648_),
    .B1(_18652_),
    .B2(_18721_),
    .X(_18722_));
 sky130_fd_sc_hd__nor2_1 _21515_ (.A(_18644_),
    .B(_18722_),
    .Y(_04002_));
 sky130_fd_sc_hd__nand2_1 _21516_ (.A(_18720_),
    .B(_18668_),
    .Y(_18723_));
 sky130_fd_sc_hd__nand2_1 _21517_ (.A(_18670_),
    .B(instr_bltu),
    .Y(_18724_));
 sky130_fd_sc_hd__a21oi_1 _21518_ (.A1(_18723_),
    .A2(_18724_),
    .B1(_18683_),
    .Y(_04001_));
 sky130_fd_sc_hd__a22o_1 _21519_ (.A1(instr_bge),
    .A2(_18687_),
    .B1(_18720_),
    .B2(_18678_),
    .X(_18725_));
 sky130_fd_sc_hd__and2_1 _21520_ (.A(_18725_),
    .B(_18333_),
    .X(_04000_));
 sky130_fd_sc_hd__a22o_1 _21521_ (.A1(instr_blt),
    .A2(_18687_),
    .B1(_18720_),
    .B2(_18688_),
    .X(_18726_));
 sky130_fd_sc_hd__and2_1 _21522_ (.A(_18726_),
    .B(_18333_),
    .X(_03999_));
 sky130_vsdinv _21523_ (.A(instr_bne),
    .Y(_18727_));
 sky130_fd_sc_hd__buf_2 _21524_ (.A(_18645_),
    .X(_18728_));
 sky130_fd_sc_hd__o2bb2a_1 _21525_ (.A1_N(_18700_),
    .A2_N(_18720_),
    .B1(_18727_),
    .B2(_18728_),
    .X(_18729_));
 sky130_fd_sc_hd__nor2_1 _21526_ (.A(_18644_),
    .B(_18729_),
    .Y(_03998_));
 sky130_fd_sc_hd__a22o_1 _21527_ (.A1(instr_beq),
    .A2(_18711_),
    .B1(_18720_),
    .B2(_18702_),
    .X(_18730_));
 sky130_fd_sc_hd__and2_1 _21528_ (.A(_18730_),
    .B(_18333_),
    .X(_03997_));
 sky130_vsdinv _21529_ (.A(\pcpi_timeout_counter[3] ),
    .Y(_18731_));
 sky130_fd_sc_hd__nor2_1 _21530_ (.A(\pcpi_timeout_counter[1] ),
    .B(\pcpi_timeout_counter[0] ),
    .Y(_18732_));
 sky130_vsdinv _21531_ (.A(_18732_),
    .Y(_18733_));
 sky130_fd_sc_hd__nor2_2 _21532_ (.A(\pcpi_timeout_counter[2] ),
    .B(_18733_),
    .Y(_18734_));
 sky130_fd_sc_hd__o21bai_1 _21533_ (.A1(_18731_),
    .A2(_18734_),
    .B1_N(_18454_),
    .Y(_03996_));
 sky130_fd_sc_hd__a21o_1 _21534_ (.A1(_18733_),
    .A2(\pcpi_timeout_counter[2] ),
    .B1(_18454_),
    .X(_18735_));
 sky130_fd_sc_hd__a21o_1 _21535_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(_18734_),
    .B1(_18735_),
    .X(_03995_));
 sky130_fd_sc_hd__o21a_1 _21536_ (.A1(\pcpi_timeout_counter[3] ),
    .A2(\pcpi_timeout_counter[2] ),
    .B1(_18732_),
    .X(_18736_));
 sky130_fd_sc_hd__a211o_1 _21537_ (.A1(\pcpi_timeout_counter[1] ),
    .A2(\pcpi_timeout_counter[0] ),
    .B1(_18454_),
    .C1(_18736_),
    .X(_03994_));
 sky130_fd_sc_hd__nand2_1 _21538_ (.A(_18734_),
    .B(_18731_),
    .Y(_18737_));
 sky130_vsdinv _21539_ (.A(\pcpi_timeout_counter[0] ),
    .Y(_18738_));
 sky130_fd_sc_hd__a21o_1 _21540_ (.A1(_18737_),
    .A2(_18738_),
    .B1(_18454_),
    .X(_03993_));
 sky130_fd_sc_hd__nor2_4 _21541_ (.A(_18312_),
    .B(_18361_),
    .Y(_00296_));
 sky130_fd_sc_hd__nor2_2 _21542_ (.A(_18630_),
    .B(_18578_),
    .Y(_18739_));
 sky130_fd_sc_hd__or4b_1 _21543_ (.A(_18478_),
    .B(_18334_),
    .C(_18552_),
    .D_N(_18739_),
    .X(_18740_));
 sky130_fd_sc_hd__a2bb2o_1 _21544_ (.A1_N(_00296_),
    .A2_N(_18740_),
    .B1(_18630_),
    .B2(_18550_),
    .X(_03992_));
 sky130_vsdinv _21545_ (.A(_00296_),
    .Y(_18741_));
 sky130_fd_sc_hd__and3_1 _21546_ (.A(_18326_),
    .B(_18330_),
    .C(\cpu_state[6] ),
    .X(_18742_));
 sky130_fd_sc_hd__a22o_1 _21547_ (.A1(mem_do_rdata),
    .A2(_18550_),
    .B1(_18741_),
    .B2(_18742_),
    .X(_03991_));
 sky130_fd_sc_hd__clkbuf_4 _21548_ (.A(_18535_),
    .X(_18743_));
 sky130_fd_sc_hd__clkbuf_2 _21549_ (.A(_18551_),
    .X(_18744_));
 sky130_fd_sc_hd__or2_1 _21550_ (.A(\reg_next_pc[31] ),
    .B(_18744_),
    .X(_18745_));
 sky130_fd_sc_hd__o211a_1 _21551_ (.A1(_02530_),
    .A2(_18743_),
    .B1(_18337_),
    .C1(_18745_),
    .X(_03990_));
 sky130_fd_sc_hd__buf_4 _21552_ (.A(_18528_),
    .X(_00322_));
 sky130_fd_sc_hd__clkbuf_2 _21553_ (.A(_18336_),
    .X(_18746_));
 sky130_fd_sc_hd__clkbuf_2 _21554_ (.A(_18551_),
    .X(_18747_));
 sky130_fd_sc_hd__or2_1 _21555_ (.A(_18747_),
    .B(\reg_next_pc[30] ),
    .X(_18748_));
 sky130_fd_sc_hd__o211a_1 _21556_ (.A1(_00322_),
    .A2(_02529_),
    .B1(_18746_),
    .C1(_18748_),
    .X(_03989_));
 sky130_fd_sc_hd__or2_1 _21557_ (.A(_18747_),
    .B(\reg_next_pc[29] ),
    .X(_18749_));
 sky130_fd_sc_hd__o211a_1 _21558_ (.A1(_00322_),
    .A2(_02527_),
    .B1(_18746_),
    .C1(_18749_),
    .X(_03988_));
 sky130_fd_sc_hd__or2_1 _21559_ (.A(_18747_),
    .B(\reg_next_pc[28] ),
    .X(_18750_));
 sky130_fd_sc_hd__o211a_1 _21560_ (.A1(_00322_),
    .A2(_02526_),
    .B1(_18746_),
    .C1(_18750_),
    .X(_03987_));
 sky130_fd_sc_hd__or2_1 _21561_ (.A(_18747_),
    .B(\reg_next_pc[27] ),
    .X(_18751_));
 sky130_fd_sc_hd__o211a_1 _21562_ (.A1(_00322_),
    .A2(_02525_),
    .B1(_18746_),
    .C1(_18751_),
    .X(_03986_));
 sky130_fd_sc_hd__or2_1 _21563_ (.A(_18747_),
    .B(\reg_next_pc[26] ),
    .X(_18752_));
 sky130_fd_sc_hd__o211a_1 _21564_ (.A1(_00322_),
    .A2(_02524_),
    .B1(_18746_),
    .C1(_18752_),
    .X(_03985_));
 sky130_fd_sc_hd__clkbuf_2 _21565_ (.A(_18528_),
    .X(_18753_));
 sky130_fd_sc_hd__buf_4 _21566_ (.A(\cpu_state[1] ),
    .X(_18754_));
 sky130_fd_sc_hd__buf_1 _21567_ (.A(_18754_),
    .X(_18755_));
 sky130_fd_sc_hd__or2_1 _21568_ (.A(_18755_),
    .B(\reg_next_pc[25] ),
    .X(_18756_));
 sky130_fd_sc_hd__o211a_1 _21569_ (.A1(_18753_),
    .A2(_02523_),
    .B1(_18746_),
    .C1(_18756_),
    .X(_03984_));
 sky130_fd_sc_hd__clkbuf_2 _21570_ (.A(_18336_),
    .X(_18757_));
 sky130_fd_sc_hd__or2_1 _21571_ (.A(_18755_),
    .B(\reg_next_pc[24] ),
    .X(_18758_));
 sky130_fd_sc_hd__o211a_1 _21572_ (.A1(_18753_),
    .A2(_02522_),
    .B1(_18757_),
    .C1(_18758_),
    .X(_03983_));
 sky130_fd_sc_hd__or2_1 _21573_ (.A(_18755_),
    .B(\reg_next_pc[23] ),
    .X(_18759_));
 sky130_fd_sc_hd__o211a_1 _21574_ (.A1(_18753_),
    .A2(_02521_),
    .B1(_18757_),
    .C1(_18759_),
    .X(_03982_));
 sky130_fd_sc_hd__or2_1 _21575_ (.A(_18755_),
    .B(\reg_next_pc[22] ),
    .X(_18760_));
 sky130_fd_sc_hd__o211a_1 _21576_ (.A1(_18753_),
    .A2(_02520_),
    .B1(_18757_),
    .C1(_18760_),
    .X(_03981_));
 sky130_fd_sc_hd__or2_1 _21577_ (.A(_18755_),
    .B(\reg_next_pc[21] ),
    .X(_18761_));
 sky130_fd_sc_hd__o211a_1 _21578_ (.A1(_18753_),
    .A2(_02519_),
    .B1(_18757_),
    .C1(_18761_),
    .X(_03980_));
 sky130_fd_sc_hd__or2_1 _21579_ (.A(_18755_),
    .B(\reg_next_pc[20] ),
    .X(_18762_));
 sky130_fd_sc_hd__o211a_1 _21580_ (.A1(_18753_),
    .A2(_02518_),
    .B1(_18757_),
    .C1(_18762_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_2 _21581_ (.A(_18528_),
    .X(_18763_));
 sky130_fd_sc_hd__buf_1 _21582_ (.A(_18551_),
    .X(_18764_));
 sky130_fd_sc_hd__or2_1 _21583_ (.A(_18764_),
    .B(\reg_next_pc[19] ),
    .X(_18765_));
 sky130_fd_sc_hd__o211a_1 _21584_ (.A1(_18763_),
    .A2(_02516_),
    .B1(_18757_),
    .C1(_18765_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_2 _21585_ (.A(_18336_),
    .X(_18766_));
 sky130_fd_sc_hd__or2_1 _21586_ (.A(_18764_),
    .B(\reg_next_pc[18] ),
    .X(_18767_));
 sky130_fd_sc_hd__o211a_1 _21587_ (.A1(_18763_),
    .A2(_02515_),
    .B1(_18766_),
    .C1(_18767_),
    .X(_03977_));
 sky130_fd_sc_hd__or2_1 _21588_ (.A(_18764_),
    .B(\reg_next_pc[17] ),
    .X(_18768_));
 sky130_fd_sc_hd__o211a_1 _21589_ (.A1(_18763_),
    .A2(_02514_),
    .B1(_18766_),
    .C1(_18768_),
    .X(_03976_));
 sky130_fd_sc_hd__or2_1 _21590_ (.A(_18764_),
    .B(\reg_next_pc[16] ),
    .X(_18769_));
 sky130_fd_sc_hd__o211a_1 _21591_ (.A1(_18763_),
    .A2(_02513_),
    .B1(_18766_),
    .C1(_18769_),
    .X(_03975_));
 sky130_fd_sc_hd__or2_1 _21592_ (.A(_18764_),
    .B(\reg_next_pc[15] ),
    .X(_18770_));
 sky130_fd_sc_hd__o211a_1 _21593_ (.A1(_18763_),
    .A2(_02512_),
    .B1(_18766_),
    .C1(_18770_),
    .X(_03974_));
 sky130_fd_sc_hd__or2_1 _21594_ (.A(_18764_),
    .B(\reg_next_pc[14] ),
    .X(_18771_));
 sky130_fd_sc_hd__o211a_1 _21595_ (.A1(_18763_),
    .A2(_02511_),
    .B1(_18766_),
    .C1(_18771_),
    .X(_03973_));
 sky130_fd_sc_hd__clkbuf_4 _21596_ (.A(_18535_),
    .X(_18772_));
 sky130_fd_sc_hd__clkbuf_2 _21597_ (.A(_18551_),
    .X(_18773_));
 sky130_fd_sc_hd__or2_1 _21598_ (.A(_18773_),
    .B(\reg_next_pc[13] ),
    .X(_18774_));
 sky130_fd_sc_hd__o211a_1 _21599_ (.A1(_18772_),
    .A2(_02510_),
    .B1(_18766_),
    .C1(_18774_),
    .X(_03972_));
 sky130_fd_sc_hd__buf_2 _21600_ (.A(_18336_),
    .X(_18775_));
 sky130_fd_sc_hd__or2_1 _21601_ (.A(_18773_),
    .B(\reg_next_pc[12] ),
    .X(_18776_));
 sky130_fd_sc_hd__o211a_1 _21602_ (.A1(_18772_),
    .A2(_02509_),
    .B1(_18775_),
    .C1(_18776_),
    .X(_03971_));
 sky130_fd_sc_hd__or2_1 _21603_ (.A(_18773_),
    .B(\reg_next_pc[11] ),
    .X(_18777_));
 sky130_fd_sc_hd__o211a_1 _21604_ (.A1(_18772_),
    .A2(_02508_),
    .B1(_18775_),
    .C1(_18777_),
    .X(_03970_));
 sky130_fd_sc_hd__or2_1 _21605_ (.A(_18773_),
    .B(\reg_next_pc[10] ),
    .X(_18778_));
 sky130_fd_sc_hd__o211a_1 _21606_ (.A1(_18772_),
    .A2(_02507_),
    .B1(_18775_),
    .C1(_18778_),
    .X(_03969_));
 sky130_fd_sc_hd__or2_1 _21607_ (.A(_18773_),
    .B(\reg_next_pc[9] ),
    .X(_18779_));
 sky130_fd_sc_hd__o211a_1 _21608_ (.A1(_18772_),
    .A2(_02537_),
    .B1(_18775_),
    .C1(_18779_),
    .X(_03968_));
 sky130_fd_sc_hd__or2_1 _21609_ (.A(_18773_),
    .B(\reg_next_pc[8] ),
    .X(_18780_));
 sky130_fd_sc_hd__o211a_1 _21610_ (.A1(_18772_),
    .A2(_02536_),
    .B1(_18775_),
    .C1(_18780_),
    .X(_03967_));
 sky130_fd_sc_hd__clkbuf_2 _21611_ (.A(_18535_),
    .X(_18781_));
 sky130_fd_sc_hd__clkbuf_2 _21612_ (.A(_18551_),
    .X(_18782_));
 sky130_fd_sc_hd__or2_1 _21613_ (.A(_18782_),
    .B(\reg_next_pc[7] ),
    .X(_18783_));
 sky130_fd_sc_hd__o211a_1 _21614_ (.A1(_18781_),
    .A2(_02535_),
    .B1(_18775_),
    .C1(_18783_),
    .X(_03966_));
 sky130_fd_sc_hd__clkbuf_4 _21615_ (.A(_18331_),
    .X(_18784_));
 sky130_fd_sc_hd__clkbuf_2 _21616_ (.A(_18784_),
    .X(_18785_));
 sky130_fd_sc_hd__or2_1 _21617_ (.A(_18782_),
    .B(\reg_next_pc[6] ),
    .X(_18786_));
 sky130_fd_sc_hd__o211a_1 _21618_ (.A1(_18781_),
    .A2(_02534_),
    .B1(_18785_),
    .C1(_18786_),
    .X(_03965_));
 sky130_fd_sc_hd__or2_1 _21619_ (.A(_18782_),
    .B(\reg_next_pc[5] ),
    .X(_18787_));
 sky130_fd_sc_hd__o211a_1 _21620_ (.A1(_18781_),
    .A2(_02533_),
    .B1(_18785_),
    .C1(_18787_),
    .X(_03964_));
 sky130_fd_sc_hd__buf_2 _21621_ (.A(_18535_),
    .X(_18788_));
 sky130_fd_sc_hd__inv_2 _21622_ (.A(\reg_next_pc[4] ),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_1 _21623_ (.A(_18788_),
    .B(_01471_),
    .Y(_18789_));
 sky130_fd_sc_hd__o211a_1 _21624_ (.A1(_18781_),
    .A2(_02532_),
    .B1(_18785_),
    .C1(_18789_),
    .X(_03963_));
 sky130_fd_sc_hd__or2_1 _21625_ (.A(_18782_),
    .B(\reg_next_pc[3] ),
    .X(_18790_));
 sky130_fd_sc_hd__o211a_1 _21626_ (.A1(_18781_),
    .A2(_02531_),
    .B1(_18785_),
    .C1(_18790_),
    .X(_03962_));
 sky130_fd_sc_hd__or2_1 _21627_ (.A(_18782_),
    .B(\reg_next_pc[2] ),
    .X(_18791_));
 sky130_fd_sc_hd__o211a_1 _21628_ (.A1(_18781_),
    .A2(_02528_),
    .B1(_18785_),
    .C1(_18791_),
    .X(_03961_));
 sky130_fd_sc_hd__or2_1 _21629_ (.A(_18782_),
    .B(\reg_next_pc[1] ),
    .X(_18792_));
 sky130_fd_sc_hd__o211a_1 _21630_ (.A1(_18743_),
    .A2(_02517_),
    .B1(_18785_),
    .C1(_18792_),
    .X(_03960_));
 sky130_fd_sc_hd__clkbuf_4 _21631_ (.A(_18744_),
    .X(_18793_));
 sky130_fd_sc_hd__clkbuf_2 _21632_ (.A(_18784_),
    .X(_18794_));
 sky130_vsdinv _21633_ (.A(_02581_),
    .Y(_18795_));
 sky130_fd_sc_hd__buf_2 _21634_ (.A(_18744_),
    .X(_18796_));
 sky130_fd_sc_hd__nand2_1 _21635_ (.A(_18795_),
    .B(_18796_),
    .Y(_18797_));
 sky130_fd_sc_hd__o211a_1 _21636_ (.A1(_18793_),
    .A2(\reg_pc[31] ),
    .B1(_18794_),
    .C1(_18797_),
    .X(_03959_));
 sky130_vsdinv _21637_ (.A(_02580_),
    .Y(_18798_));
 sky130_fd_sc_hd__clkbuf_2 _21638_ (.A(_18754_),
    .X(_18799_));
 sky130_fd_sc_hd__nand2_1 _21639_ (.A(_18798_),
    .B(_18799_),
    .Y(_18800_));
 sky130_fd_sc_hd__o211a_1 _21640_ (.A1(_18793_),
    .A2(\reg_pc[30] ),
    .B1(_18794_),
    .C1(_18800_),
    .X(_03958_));
 sky130_vsdinv _21641_ (.A(_02579_),
    .Y(_18801_));
 sky130_fd_sc_hd__nand2_1 _21642_ (.A(_18801_),
    .B(_18799_),
    .Y(_18802_));
 sky130_fd_sc_hd__o211a_1 _21643_ (.A1(_18793_),
    .A2(\reg_pc[29] ),
    .B1(_18794_),
    .C1(_18802_),
    .X(_03957_));
 sky130_vsdinv _21644_ (.A(_02578_),
    .Y(_18803_));
 sky130_fd_sc_hd__nand2_1 _21645_ (.A(_18803_),
    .B(_18799_),
    .Y(_18804_));
 sky130_fd_sc_hd__o211a_1 _21646_ (.A1(_18793_),
    .A2(\reg_pc[28] ),
    .B1(_18794_),
    .C1(_18804_),
    .X(_03956_));
 sky130_vsdinv _21647_ (.A(_02577_),
    .Y(_18805_));
 sky130_fd_sc_hd__nand2_1 _21648_ (.A(_18805_),
    .B(_18799_),
    .Y(_18806_));
 sky130_fd_sc_hd__o211a_1 _21649_ (.A1(_18793_),
    .A2(\reg_pc[27] ),
    .B1(_18794_),
    .C1(_18806_),
    .X(_03955_));
 sky130_fd_sc_hd__clkbuf_2 _21650_ (.A(_18744_),
    .X(_18807_));
 sky130_vsdinv _21651_ (.A(_02576_),
    .Y(_18808_));
 sky130_fd_sc_hd__nand2_1 _21652_ (.A(_18808_),
    .B(_18799_),
    .Y(_18809_));
 sky130_fd_sc_hd__o211a_1 _21653_ (.A1(_18807_),
    .A2(\reg_pc[26] ),
    .B1(_18794_),
    .C1(_18809_),
    .X(_03954_));
 sky130_fd_sc_hd__clkbuf_2 _21654_ (.A(_18784_),
    .X(_18810_));
 sky130_vsdinv _21655_ (.A(_02575_),
    .Y(_18811_));
 sky130_fd_sc_hd__nand2_1 _21656_ (.A(_18811_),
    .B(_18799_),
    .Y(_18812_));
 sky130_fd_sc_hd__o211a_1 _21657_ (.A1(_18807_),
    .A2(\reg_pc[25] ),
    .B1(_18810_),
    .C1(_18812_),
    .X(_03953_));
 sky130_vsdinv _21658_ (.A(_02574_),
    .Y(_18813_));
 sky130_fd_sc_hd__clkbuf_2 _21659_ (.A(_18754_),
    .X(_18814_));
 sky130_fd_sc_hd__nand2_1 _21660_ (.A(_18813_),
    .B(_18814_),
    .Y(_18815_));
 sky130_fd_sc_hd__o211a_1 _21661_ (.A1(_18807_),
    .A2(\reg_pc[24] ),
    .B1(_18810_),
    .C1(_18815_),
    .X(_03952_));
 sky130_vsdinv _21662_ (.A(_02573_),
    .Y(_18816_));
 sky130_fd_sc_hd__nand2_1 _21663_ (.A(_18816_),
    .B(_18814_),
    .Y(_18817_));
 sky130_fd_sc_hd__o211a_1 _21664_ (.A1(_18807_),
    .A2(\reg_pc[23] ),
    .B1(_18810_),
    .C1(_18817_),
    .X(_03951_));
 sky130_vsdinv _21665_ (.A(_02572_),
    .Y(_18818_));
 sky130_fd_sc_hd__nand2_1 _21666_ (.A(_18818_),
    .B(_18814_),
    .Y(_18819_));
 sky130_fd_sc_hd__o211a_1 _21667_ (.A1(_18807_),
    .A2(\reg_pc[22] ),
    .B1(_18810_),
    .C1(_18819_),
    .X(_03950_));
 sky130_vsdinv _21668_ (.A(_02570_),
    .Y(_18820_));
 sky130_fd_sc_hd__nand2_1 _21669_ (.A(_18820_),
    .B(_18814_),
    .Y(_18821_));
 sky130_fd_sc_hd__o211a_1 _21670_ (.A1(_18807_),
    .A2(\reg_pc[21] ),
    .B1(_18810_),
    .C1(_18821_),
    .X(_03949_));
 sky130_fd_sc_hd__buf_2 _21671_ (.A(_18744_),
    .X(_18822_));
 sky130_vsdinv _21672_ (.A(_02569_),
    .Y(_18823_));
 sky130_fd_sc_hd__nand2_1 _21673_ (.A(_18823_),
    .B(_18814_),
    .Y(_18824_));
 sky130_fd_sc_hd__o211a_1 _21674_ (.A1(_18822_),
    .A2(\reg_pc[20] ),
    .B1(_18810_),
    .C1(_18824_),
    .X(_03948_));
 sky130_fd_sc_hd__clkbuf_2 _21675_ (.A(_18784_),
    .X(_18825_));
 sky130_vsdinv _21676_ (.A(_02568_),
    .Y(_18826_));
 sky130_fd_sc_hd__nand2_1 _21677_ (.A(_18826_),
    .B(_18814_),
    .Y(_18827_));
 sky130_fd_sc_hd__o211a_1 _21678_ (.A1(_18822_),
    .A2(\reg_pc[19] ),
    .B1(_18825_),
    .C1(_18827_),
    .X(_03947_));
 sky130_vsdinv _21679_ (.A(_02567_),
    .Y(_18828_));
 sky130_fd_sc_hd__clkbuf_2 _21680_ (.A(_18754_),
    .X(_18829_));
 sky130_fd_sc_hd__nand2_1 _21681_ (.A(_18828_),
    .B(_18829_),
    .Y(_18830_));
 sky130_fd_sc_hd__o211a_1 _21682_ (.A1(_18822_),
    .A2(\reg_pc[18] ),
    .B1(_18825_),
    .C1(_18830_),
    .X(_03946_));
 sky130_vsdinv _21683_ (.A(_02566_),
    .Y(_18831_));
 sky130_fd_sc_hd__nand2_1 _21684_ (.A(_18831_),
    .B(_18829_),
    .Y(_18832_));
 sky130_fd_sc_hd__o211a_1 _21685_ (.A1(_18822_),
    .A2(\reg_pc[17] ),
    .B1(_18825_),
    .C1(_18832_),
    .X(_03945_));
 sky130_vsdinv _21686_ (.A(_02565_),
    .Y(_18833_));
 sky130_fd_sc_hd__nand2_1 _21687_ (.A(_18833_),
    .B(_18829_),
    .Y(_18834_));
 sky130_fd_sc_hd__o211a_1 _21688_ (.A1(_18822_),
    .A2(\reg_pc[16] ),
    .B1(_18825_),
    .C1(_18834_),
    .X(_03944_));
 sky130_vsdinv _21689_ (.A(_02564_),
    .Y(_18835_));
 sky130_fd_sc_hd__nand2_1 _21690_ (.A(_18835_),
    .B(_18829_),
    .Y(_18836_));
 sky130_fd_sc_hd__o211a_1 _21691_ (.A1(_18822_),
    .A2(\reg_pc[15] ),
    .B1(_18825_),
    .C1(_18836_),
    .X(_03943_));
 sky130_fd_sc_hd__buf_2 _21692_ (.A(_18744_),
    .X(_18837_));
 sky130_vsdinv _21693_ (.A(_02563_),
    .Y(_18838_));
 sky130_fd_sc_hd__nand2_1 _21694_ (.A(_18838_),
    .B(_18829_),
    .Y(_18839_));
 sky130_fd_sc_hd__o211a_1 _21695_ (.A1(_18837_),
    .A2(\reg_pc[14] ),
    .B1(_18825_),
    .C1(_18839_),
    .X(_03942_));
 sky130_fd_sc_hd__buf_2 _21696_ (.A(_18784_),
    .X(_18840_));
 sky130_vsdinv _21697_ (.A(_02562_),
    .Y(_18841_));
 sky130_fd_sc_hd__nand2_1 _21698_ (.A(_18841_),
    .B(_18829_),
    .Y(_18842_));
 sky130_fd_sc_hd__o211a_1 _21699_ (.A1(_18837_),
    .A2(\reg_pc[13] ),
    .B1(_18840_),
    .C1(_18842_),
    .X(_03941_));
 sky130_vsdinv _21700_ (.A(_02561_),
    .Y(_18843_));
 sky130_fd_sc_hd__buf_2 _21701_ (.A(_18754_),
    .X(_18844_));
 sky130_fd_sc_hd__nand2_1 _21702_ (.A(_18843_),
    .B(_18844_),
    .Y(_18845_));
 sky130_fd_sc_hd__o211a_1 _21703_ (.A1(_18837_),
    .A2(\reg_pc[12] ),
    .B1(_18840_),
    .C1(_18845_),
    .X(_03940_));
 sky130_vsdinv _21704_ (.A(_02589_),
    .Y(_18846_));
 sky130_fd_sc_hd__nand2_1 _21705_ (.A(_18846_),
    .B(_18844_),
    .Y(_18847_));
 sky130_fd_sc_hd__o211a_1 _21706_ (.A1(_18837_),
    .A2(\reg_pc[11] ),
    .B1(_18840_),
    .C1(_18847_),
    .X(_03939_));
 sky130_vsdinv _21707_ (.A(_02588_),
    .Y(_18848_));
 sky130_fd_sc_hd__nand2_1 _21708_ (.A(_18848_),
    .B(_18844_),
    .Y(_18849_));
 sky130_fd_sc_hd__o211a_1 _21709_ (.A1(_18837_),
    .A2(\reg_pc[10] ),
    .B1(_18840_),
    .C1(_18849_),
    .X(_03938_));
 sky130_vsdinv _21710_ (.A(\reg_pc[9] ),
    .Y(_18850_));
 sky130_fd_sc_hd__nand2_1 _21711_ (.A(_18788_),
    .B(_18850_),
    .Y(_18851_));
 sky130_fd_sc_hd__o211a_1 _21712_ (.A1(_18743_),
    .A2(_02587_),
    .B1(_18840_),
    .C1(_18851_),
    .X(_03937_));
 sky130_vsdinv _21713_ (.A(_02586_),
    .Y(_18852_));
 sky130_fd_sc_hd__nand2_1 _21714_ (.A(_18852_),
    .B(_18844_),
    .Y(_18853_));
 sky130_fd_sc_hd__o211a_1 _21715_ (.A1(_18837_),
    .A2(\reg_pc[8] ),
    .B1(_18840_),
    .C1(_18853_),
    .X(_03936_));
 sky130_fd_sc_hd__clkbuf_2 _21716_ (.A(_18784_),
    .X(_18854_));
 sky130_vsdinv _21717_ (.A(\reg_pc[7] ),
    .Y(_18855_));
 sky130_fd_sc_hd__nand2_1 _21718_ (.A(_18788_),
    .B(_18855_),
    .Y(_18856_));
 sky130_fd_sc_hd__o211a_1 _21719_ (.A1(_18743_),
    .A2(_02585_),
    .B1(_18854_),
    .C1(_18856_),
    .X(_03935_));
 sky130_vsdinv _21720_ (.A(_02584_),
    .Y(_18857_));
 sky130_fd_sc_hd__nand2_1 _21721_ (.A(_18857_),
    .B(_18844_),
    .Y(_18858_));
 sky130_fd_sc_hd__o211a_1 _21722_ (.A1(_18796_),
    .A2(\reg_pc[6] ),
    .B1(_18854_),
    .C1(_18858_),
    .X(_03934_));
 sky130_vsdinv _21723_ (.A(\reg_pc[5] ),
    .Y(_18859_));
 sky130_fd_sc_hd__nand2_1 _21724_ (.A(_18788_),
    .B(_18859_),
    .Y(_18860_));
 sky130_fd_sc_hd__o211a_1 _21725_ (.A1(_18743_),
    .A2(_02583_),
    .B1(_18854_),
    .C1(_18860_),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_1 _21726_ (.A(_18796_),
    .B(_01475_),
    .Y(_18861_));
 sky130_fd_sc_hd__o211a_1 _21727_ (.A1(_18796_),
    .A2(\reg_pc[4] ),
    .B1(_18854_),
    .C1(_18861_),
    .X(_03932_));
 sky130_fd_sc_hd__inv_2 _21728_ (.A(_01475_),
    .Y(_02582_));
 sky130_vsdinv _21729_ (.A(_02571_),
    .Y(_18862_));
 sky130_fd_sc_hd__nand2_1 _21730_ (.A(_18862_),
    .B(_18844_),
    .Y(_18863_));
 sky130_fd_sc_hd__o211a_1 _21731_ (.A1(_18796_),
    .A2(\reg_pc[3] ),
    .B1(_18854_),
    .C1(_18863_),
    .X(_03931_));
 sky130_fd_sc_hd__inv_2 _21732_ (.A(_02560_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_1 _21733_ (.A(_01561_),
    .B(_18747_),
    .Y(_18864_));
 sky130_fd_sc_hd__o211a_1 _21734_ (.A1(_18796_),
    .A2(\reg_pc[2] ),
    .B1(_18854_),
    .C1(_18864_),
    .X(_03930_));
 sky130_fd_sc_hd__clkbuf_2 _21735_ (.A(_18331_),
    .X(_18865_));
 sky130_fd_sc_hd__buf_4 _21736_ (.A(_18865_),
    .X(_18866_));
 sky130_vsdinv _21737_ (.A(\reg_pc[1] ),
    .Y(_18867_));
 sky130_fd_sc_hd__nand2_1 _21738_ (.A(_18788_),
    .B(_18867_),
    .Y(_18868_));
 sky130_fd_sc_hd__o211a_1 _21739_ (.A1(_18743_),
    .A2(_02590_),
    .B1(_18866_),
    .C1(_18868_),
    .X(_03929_));
 sky130_fd_sc_hd__clkbuf_2 _21740_ (.A(_18532_),
    .X(_18869_));
 sky130_fd_sc_hd__clkbuf_4 _21741_ (.A(_18869_),
    .X(_18870_));
 sky130_vsdinv _21742_ (.A(\count_instr[58] ),
    .Y(_18871_));
 sky130_fd_sc_hd__nand2_1 _21743_ (.A(\count_instr[57] ),
    .B(\count_instr[56] ),
    .Y(_18872_));
 sky130_fd_sc_hd__nand2_1 _21744_ (.A(\count_instr[47] ),
    .B(\count_instr[46] ),
    .Y(_18873_));
 sky130_vsdinv _21745_ (.A(\count_instr[48] ),
    .Y(_18874_));
 sky130_vsdinv _21746_ (.A(\count_instr[45] ),
    .Y(_18875_));
 sky130_vsdinv _21747_ (.A(\count_instr[44] ),
    .Y(_18876_));
 sky130_fd_sc_hd__or4_4 _21748_ (.A(_18873_),
    .B(_18874_),
    .C(_18875_),
    .D(_18876_),
    .X(_18877_));
 sky130_fd_sc_hd__nand2_1 _21749_ (.A(\count_instr[50] ),
    .B(\count_instr[49] ),
    .Y(_18878_));
 sky130_fd_sc_hd__and2_1 _21750_ (.A(\count_instr[36] ),
    .B(\count_instr[35] ),
    .X(_18879_));
 sky130_vsdinv _21751_ (.A(_18879_),
    .Y(_18880_));
 sky130_fd_sc_hd__and3_1 _21752_ (.A(\count_instr[39] ),
    .B(\count_instr[38] ),
    .C(\count_instr[37] ),
    .X(_18881_));
 sky130_vsdinv _21753_ (.A(_18881_),
    .Y(_18882_));
 sky130_vsdinv _21754_ (.A(\count_instr[26] ),
    .Y(_18883_));
 sky130_vsdinv _21755_ (.A(\count_instr[25] ),
    .Y(_18884_));
 sky130_fd_sc_hd__nor2_1 _21756_ (.A(_18883_),
    .B(_18884_),
    .Y(_18885_));
 sky130_vsdinv _21757_ (.A(_18885_),
    .Y(_18886_));
 sky130_fd_sc_hd__and3_1 _21758_ (.A(\count_instr[31] ),
    .B(\count_instr[30] ),
    .C(\count_instr[29] ),
    .X(_18887_));
 sky130_fd_sc_hd__and3_1 _21759_ (.A(_18887_),
    .B(\count_instr[28] ),
    .C(\count_instr[27] ),
    .X(_18888_));
 sky130_vsdinv _21760_ (.A(_18888_),
    .Y(_18889_));
 sky130_vsdinv _21761_ (.A(\count_instr[13] ),
    .Y(_18890_));
 sky130_fd_sc_hd__and4_1 _21762_ (.A(\count_instr[12] ),
    .B(\count_instr[11] ),
    .C(\count_instr[10] ),
    .D(\count_instr[9] ),
    .X(_18891_));
 sky130_fd_sc_hd__and3_1 _21763_ (.A(\count_instr[4] ),
    .B(\count_instr[3] ),
    .C(\count_instr[0] ),
    .X(_18892_));
 sky130_fd_sc_hd__and4_1 _21764_ (.A(_18891_),
    .B(\count_instr[2] ),
    .C(_18892_),
    .D(\count_instr[1] ),
    .X(_18893_));
 sky130_fd_sc_hd__and3_1 _21765_ (.A(\count_instr[8] ),
    .B(\count_instr[7] ),
    .C(\count_instr[6] ),
    .X(_18894_));
 sky130_fd_sc_hd__and3_1 _21766_ (.A(_18893_),
    .B(\count_instr[5] ),
    .C(_18894_),
    .X(_18895_));
 sky130_fd_sc_hd__nand2_2 _21767_ (.A(_18448_),
    .B(_18895_),
    .Y(_18896_));
 sky130_fd_sc_hd__nor2_2 _21768_ (.A(_18890_),
    .B(_18896_),
    .Y(_18897_));
 sky130_fd_sc_hd__and3_1 _21769_ (.A(_18897_),
    .B(\count_instr[15] ),
    .C(\count_instr[14] ),
    .X(_18898_));
 sky130_fd_sc_hd__and4_1 _21770_ (.A(_18898_),
    .B(\count_instr[18] ),
    .C(\count_instr[17] ),
    .D(\count_instr[16] ),
    .X(_18899_));
 sky130_vsdinv _21771_ (.A(\count_instr[20] ),
    .Y(_18900_));
 sky130_vsdinv _21772_ (.A(\count_instr[19] ),
    .Y(_18901_));
 sky130_fd_sc_hd__nor2_1 _21773_ (.A(_18900_),
    .B(_18901_),
    .Y(_18902_));
 sky130_fd_sc_hd__and3_2 _21774_ (.A(_18899_),
    .B(\count_instr[21] ),
    .C(_18902_),
    .X(_18903_));
 sky130_vsdinv _21775_ (.A(\count_instr[23] ),
    .Y(_18904_));
 sky130_vsdinv _21776_ (.A(\count_instr[22] ),
    .Y(_18905_));
 sky130_fd_sc_hd__nor2_2 _21777_ (.A(_18904_),
    .B(_18905_),
    .Y(_18906_));
 sky130_fd_sc_hd__nand3_4 _21778_ (.A(_18903_),
    .B(\count_instr[24] ),
    .C(_18906_),
    .Y(_18907_));
 sky130_fd_sc_hd__nor3_4 _21779_ (.A(_18886_),
    .B(_18889_),
    .C(_18907_),
    .Y(_18908_));
 sky130_vsdinv _21780_ (.A(\count_instr[34] ),
    .Y(_18909_));
 sky130_vsdinv _21781_ (.A(\count_instr[33] ),
    .Y(_18910_));
 sky130_fd_sc_hd__nor2_2 _21782_ (.A(_18909_),
    .B(_18910_),
    .Y(_18911_));
 sky130_fd_sc_hd__nand3_4 _21783_ (.A(_18908_),
    .B(\count_instr[32] ),
    .C(_18911_),
    .Y(_18912_));
 sky130_fd_sc_hd__nor3_4 _21784_ (.A(_18880_),
    .B(_18882_),
    .C(_18912_),
    .Y(_18913_));
 sky130_vsdinv _21785_ (.A(\count_instr[41] ),
    .Y(_18914_));
 sky130_vsdinv _21786_ (.A(\count_instr[40] ),
    .Y(_18915_));
 sky130_fd_sc_hd__nor2_2 _21787_ (.A(_18914_),
    .B(_18915_),
    .Y(_18916_));
 sky130_fd_sc_hd__and2_1 _21788_ (.A(\count_instr[43] ),
    .B(\count_instr[42] ),
    .X(_18917_));
 sky130_fd_sc_hd__nand3_4 _21789_ (.A(_18913_),
    .B(_18916_),
    .C(_18917_),
    .Y(_18918_));
 sky130_fd_sc_hd__nor3_4 _21790_ (.A(_18877_),
    .B(_18878_),
    .C(_18918_),
    .Y(_18919_));
 sky130_vsdinv _21791_ (.A(\count_instr[52] ),
    .Y(_18920_));
 sky130_vsdinv _21792_ (.A(\count_instr[51] ),
    .Y(_18921_));
 sky130_fd_sc_hd__nor2_2 _21793_ (.A(_18920_),
    .B(_18921_),
    .Y(_18922_));
 sky130_fd_sc_hd__and3_1 _21794_ (.A(\count_instr[55] ),
    .B(\count_instr[54] ),
    .C(\count_instr[53] ),
    .X(_18923_));
 sky130_fd_sc_hd__nand3_4 _21795_ (.A(_18919_),
    .B(_18922_),
    .C(_18923_),
    .Y(_18924_));
 sky130_fd_sc_hd__nor3_4 _21796_ (.A(_18871_),
    .B(_18872_),
    .C(_18924_),
    .Y(_18925_));
 sky130_fd_sc_hd__clkbuf_2 _21797_ (.A(_18925_),
    .X(_18926_));
 sky130_fd_sc_hd__clkbuf_2 _21798_ (.A(\count_instr[59] ),
    .X(_18927_));
 sky130_fd_sc_hd__and2_1 _21799_ (.A(\count_instr[61] ),
    .B(\count_instr[60] ),
    .X(_18928_));
 sky130_fd_sc_hd__a41oi_1 _21800_ (.A1(\count_instr[62] ),
    .A2(_18926_),
    .A3(_18927_),
    .A4(_18928_),
    .B1(\count_instr[63] ),
    .Y(_18929_));
 sky130_vsdinv _21801_ (.A(\count_instr[63] ),
    .Y(_18930_));
 sky130_vsdinv _21802_ (.A(\count_instr[62] ),
    .Y(_18931_));
 sky130_fd_sc_hd__nand3_4 _21803_ (.A(_18925_),
    .B(\count_instr[59] ),
    .C(_18928_),
    .Y(_18932_));
 sky130_fd_sc_hd__nor3_1 _21804_ (.A(_18930_),
    .B(_18931_),
    .C(_18932_),
    .Y(_18933_));
 sky130_fd_sc_hd__nor3_1 _21805_ (.A(_18870_),
    .B(_18929_),
    .C(_18933_),
    .Y(_03928_));
 sky130_fd_sc_hd__buf_2 _21806_ (.A(_18330_),
    .X(_18934_));
 sky130_fd_sc_hd__clkbuf_2 _21807_ (.A(_18934_),
    .X(_18935_));
 sky130_fd_sc_hd__o21ai_1 _21808_ (.A1(_18931_),
    .A2(_18932_),
    .B1(_18935_),
    .Y(_18936_));
 sky130_fd_sc_hd__a21oi_1 _21809_ (.A1(_18931_),
    .A2(_18932_),
    .B1(_18936_),
    .Y(_03927_));
 sky130_fd_sc_hd__a31o_1 _21810_ (.A1(_18926_),
    .A2(\count_instr[60] ),
    .A3(_18927_),
    .B1(\count_instr[61] ),
    .X(_18937_));
 sky130_fd_sc_hd__buf_4 _21811_ (.A(_18332_),
    .X(_18938_));
 sky130_fd_sc_hd__and3_1 _21812_ (.A(_18937_),
    .B(_18938_),
    .C(_18932_),
    .X(_03926_));
 sky130_vsdinv _21813_ (.A(\count_instr[60] ),
    .Y(_18939_));
 sky130_fd_sc_hd__nand2_1 _21814_ (.A(_18926_),
    .B(_18927_),
    .Y(_18940_));
 sky130_fd_sc_hd__a31o_1 _21815_ (.A1(_18926_),
    .A2(\count_instr[60] ),
    .A3(_18927_),
    .B1(_18869_),
    .X(_18941_));
 sky130_fd_sc_hd__a21oi_1 _21816_ (.A1(_18939_),
    .A2(_18940_),
    .B1(_18941_),
    .Y(_03925_));
 sky130_fd_sc_hd__or2_1 _21817_ (.A(_18927_),
    .B(_18926_),
    .X(_18942_));
 sky130_fd_sc_hd__clkbuf_2 _21818_ (.A(_18332_),
    .X(_18943_));
 sky130_fd_sc_hd__and3_1 _21819_ (.A(_18942_),
    .B(_18943_),
    .C(_18940_),
    .X(_03924_));
 sky130_vsdinv _21820_ (.A(\count_instr[56] ),
    .Y(_18944_));
 sky130_fd_sc_hd__nor2_1 _21821_ (.A(_18944_),
    .B(_18924_),
    .Y(_18945_));
 sky130_fd_sc_hd__nand2_1 _21822_ (.A(_18945_),
    .B(\count_instr[57] ),
    .Y(_18946_));
 sky130_fd_sc_hd__or2_1 _21823_ (.A(_18869_),
    .B(_18926_),
    .X(_18947_));
 sky130_fd_sc_hd__a21oi_1 _21824_ (.A1(_18871_),
    .A2(_18946_),
    .B1(_18947_),
    .Y(_03923_));
 sky130_fd_sc_hd__or2_1 _21825_ (.A(\count_instr[57] ),
    .B(_18945_),
    .X(_18948_));
 sky130_fd_sc_hd__and3_1 _21826_ (.A(_18948_),
    .B(_18943_),
    .C(_18946_),
    .X(_03922_));
 sky130_fd_sc_hd__or2_1 _21827_ (.A(_18869_),
    .B(_18945_),
    .X(_18949_));
 sky130_fd_sc_hd__a21oi_1 _21828_ (.A1(_18944_),
    .A2(_18924_),
    .B1(_18949_),
    .Y(_03921_));
 sky130_vsdinv _21829_ (.A(\count_instr[54] ),
    .Y(_18950_));
 sky130_fd_sc_hd__and2_1 _21830_ (.A(_18919_),
    .B(_18922_),
    .X(_18951_));
 sky130_fd_sc_hd__nand2_1 _21831_ (.A(_18951_),
    .B(\count_instr[53] ),
    .Y(_18952_));
 sky130_fd_sc_hd__or2_1 _21832_ (.A(_18950_),
    .B(_18952_),
    .X(_18953_));
 sky130_vsdinv _21833_ (.A(\count_instr[55] ),
    .Y(_18954_));
 sky130_fd_sc_hd__nand2_1 _21834_ (.A(_18924_),
    .B(_18695_),
    .Y(_18955_));
 sky130_fd_sc_hd__a21oi_1 _21835_ (.A1(_18953_),
    .A2(_18954_),
    .B1(_18955_),
    .Y(_03920_));
 sky130_fd_sc_hd__nand2_1 _21836_ (.A(_18952_),
    .B(_18950_),
    .Y(_18956_));
 sky130_fd_sc_hd__and3_1 _21837_ (.A(_18953_),
    .B(_18943_),
    .C(_18956_),
    .X(_03919_));
 sky130_fd_sc_hd__or2_1 _21838_ (.A(\count_instr[53] ),
    .B(_18951_),
    .X(_18957_));
 sky130_fd_sc_hd__and3_1 _21839_ (.A(_18957_),
    .B(_18943_),
    .C(_18952_),
    .X(_03918_));
 sky130_vsdinv _21840_ (.A(_18919_),
    .Y(_18958_));
 sky130_fd_sc_hd__nor2_1 _21841_ (.A(_18921_),
    .B(_18958_),
    .Y(_18959_));
 sky130_vsdinv _21842_ (.A(_18951_),
    .Y(_18960_));
 sky130_fd_sc_hd__o211a_1 _21843_ (.A1(\count_instr[52] ),
    .A2(_18959_),
    .B1(_18866_),
    .C1(_18960_),
    .X(_03917_));
 sky130_fd_sc_hd__nor2_1 _21844_ (.A(_18598_),
    .B(_18959_),
    .Y(_18961_));
 sky130_fd_sc_hd__o21a_1 _21845_ (.A1(\count_instr[51] ),
    .A2(_18919_),
    .B1(_18961_),
    .X(_03916_));
 sky130_fd_sc_hd__nor2_1 _21846_ (.A(_18877_),
    .B(_18918_),
    .Y(_18962_));
 sky130_fd_sc_hd__nand2_1 _21847_ (.A(_18962_),
    .B(\count_instr[49] ),
    .Y(_18963_));
 sky130_vsdinv _21848_ (.A(\count_instr[50] ),
    .Y(_18964_));
 sky130_fd_sc_hd__nand2_1 _21849_ (.A(_18963_),
    .B(_18964_),
    .Y(_18965_));
 sky130_fd_sc_hd__and3_1 _21850_ (.A(_18965_),
    .B(_18943_),
    .C(_18958_),
    .X(_03915_));
 sky130_fd_sc_hd__or2_1 _21851_ (.A(\count_instr[49] ),
    .B(_18962_),
    .X(_18966_));
 sky130_fd_sc_hd__and3_1 _21852_ (.A(_18966_),
    .B(_18943_),
    .C(_18963_),
    .X(_03914_));
 sky130_vsdinv _21853_ (.A(\count_instr[47] ),
    .Y(_18967_));
 sky130_vsdinv _21854_ (.A(\count_instr[46] ),
    .Y(_18968_));
 sky130_fd_sc_hd__or4_4 _21855_ (.A(_18968_),
    .B(_18875_),
    .C(_18876_),
    .D(_18918_),
    .X(_18969_));
 sky130_fd_sc_hd__or2_1 _21856_ (.A(_18967_),
    .B(_18969_),
    .X(_18970_));
 sky130_fd_sc_hd__a211oi_1 _21857_ (.A1(_18970_),
    .A2(_18874_),
    .B1(_18870_),
    .C1(_18962_),
    .Y(_03913_));
 sky130_fd_sc_hd__buf_1 _21858_ (.A(_18332_),
    .X(_18971_));
 sky130_fd_sc_hd__nand2_1 _21859_ (.A(_18969_),
    .B(_18967_),
    .Y(_18972_));
 sky130_fd_sc_hd__and3_1 _21860_ (.A(_18970_),
    .B(_18971_),
    .C(_18972_),
    .X(_03912_));
 sky130_fd_sc_hd__or2_1 _21861_ (.A(_18876_),
    .B(_18918_),
    .X(_18973_));
 sky130_fd_sc_hd__or2_1 _21862_ (.A(_18875_),
    .B(_18973_),
    .X(_18974_));
 sky130_fd_sc_hd__nand2_1 _21863_ (.A(_18974_),
    .B(_18968_),
    .Y(_18975_));
 sky130_fd_sc_hd__and3_1 _21864_ (.A(_18975_),
    .B(_18971_),
    .C(_18969_),
    .X(_03911_));
 sky130_fd_sc_hd__nand2_1 _21865_ (.A(_18973_),
    .B(_18875_),
    .Y(_18976_));
 sky130_fd_sc_hd__and3_1 _21866_ (.A(_18974_),
    .B(_18971_),
    .C(_18976_),
    .X(_03910_));
 sky130_fd_sc_hd__nand2_1 _21867_ (.A(_18918_),
    .B(_18876_),
    .Y(_18977_));
 sky130_fd_sc_hd__and3_1 _21868_ (.A(_18973_),
    .B(_18971_),
    .C(_18977_),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_1 _21869_ (.A(_18913_),
    .B(\count_instr[40] ),
    .Y(_18978_));
 sky130_fd_sc_hd__nor2_1 _21870_ (.A(_18914_),
    .B(_18978_),
    .Y(_18979_));
 sky130_fd_sc_hd__nand2_1 _21871_ (.A(_18979_),
    .B(\count_instr[42] ),
    .Y(_18980_));
 sky130_vsdinv _21872_ (.A(\count_instr[43] ),
    .Y(_18981_));
 sky130_fd_sc_hd__nand2_1 _21873_ (.A(_18980_),
    .B(_18981_),
    .Y(_18982_));
 sky130_fd_sc_hd__and3_1 _21874_ (.A(_18982_),
    .B(_18971_),
    .C(_18918_),
    .X(_03908_));
 sky130_fd_sc_hd__or2_1 _21875_ (.A(\count_instr[42] ),
    .B(_18979_),
    .X(_18983_));
 sky130_fd_sc_hd__and3_1 _21876_ (.A(_18983_),
    .B(_18971_),
    .C(_18980_),
    .X(_03907_));
 sky130_fd_sc_hd__buf_2 _21877_ (.A(_18578_),
    .X(_18984_));
 sky130_fd_sc_hd__or2_1 _21878_ (.A(_18984_),
    .B(_18979_),
    .X(_18985_));
 sky130_fd_sc_hd__a21oi_1 _21879_ (.A1(_18914_),
    .A2(_18978_),
    .B1(_18985_),
    .Y(_03906_));
 sky130_vsdinv _21880_ (.A(_18913_),
    .Y(_18986_));
 sky130_fd_sc_hd__nand2_1 _21881_ (.A(_18986_),
    .B(_18915_),
    .Y(_18987_));
 sky130_fd_sc_hd__clkbuf_2 _21882_ (.A(_18332_),
    .X(_18988_));
 sky130_fd_sc_hd__and3_1 _21883_ (.A(_18987_),
    .B(_18988_),
    .C(_18978_),
    .X(_03905_));
 sky130_vsdinv _21884_ (.A(\count_instr[38] ),
    .Y(_18989_));
 sky130_fd_sc_hd__nor2_1 _21885_ (.A(_18880_),
    .B(_18912_),
    .Y(_18990_));
 sky130_fd_sc_hd__nand2_1 _21886_ (.A(_18990_),
    .B(\count_instr[37] ),
    .Y(_18991_));
 sky130_fd_sc_hd__nor2_1 _21887_ (.A(_18989_),
    .B(_18991_),
    .Y(_18992_));
 sky130_fd_sc_hd__o211a_1 _21888_ (.A1(\count_instr[39] ),
    .A2(_18992_),
    .B1(_18866_),
    .C1(_18986_),
    .X(_03904_));
 sky130_fd_sc_hd__or2_1 _21889_ (.A(_18984_),
    .B(_18992_),
    .X(_18993_));
 sky130_fd_sc_hd__a21oi_1 _21890_ (.A1(_18989_),
    .A2(_18991_),
    .B1(_18993_),
    .Y(_03903_));
 sky130_vsdinv _21891_ (.A(_18990_),
    .Y(_18994_));
 sky130_vsdinv _21892_ (.A(\count_instr[37] ),
    .Y(_18995_));
 sky130_fd_sc_hd__nand2_1 _21893_ (.A(_18994_),
    .B(_18995_),
    .Y(_18996_));
 sky130_fd_sc_hd__and3_1 _21894_ (.A(_18996_),
    .B(_18988_),
    .C(_18991_),
    .X(_03902_));
 sky130_vsdinv _21895_ (.A(\count_instr[35] ),
    .Y(_18997_));
 sky130_fd_sc_hd__nor2_1 _21896_ (.A(_18997_),
    .B(_18912_),
    .Y(_18998_));
 sky130_fd_sc_hd__o211a_1 _21897_ (.A1(\count_instr[36] ),
    .A2(_18998_),
    .B1(_18866_),
    .C1(_18994_),
    .X(_03901_));
 sky130_fd_sc_hd__or2_1 _21898_ (.A(_18984_),
    .B(_18998_),
    .X(_18999_));
 sky130_fd_sc_hd__a21oi_1 _21899_ (.A1(_18997_),
    .A2(_18912_),
    .B1(_18999_),
    .Y(_03900_));
 sky130_vsdinv _21900_ (.A(\count_instr[32] ),
    .Y(_19000_));
 sky130_vsdinv _21901_ (.A(_18908_),
    .Y(_19001_));
 sky130_fd_sc_hd__nor2_1 _21902_ (.A(_19000_),
    .B(_19001_),
    .Y(_19002_));
 sky130_fd_sc_hd__nand2_1 _21903_ (.A(_19002_),
    .B(\count_instr[33] ),
    .Y(_19003_));
 sky130_fd_sc_hd__nand2_1 _21904_ (.A(_19003_),
    .B(_18909_),
    .Y(_19004_));
 sky130_fd_sc_hd__and3_1 _21905_ (.A(_19004_),
    .B(_18988_),
    .C(_18912_),
    .X(_03899_));
 sky130_vsdinv _21906_ (.A(_19002_),
    .Y(_19005_));
 sky130_fd_sc_hd__nand2_1 _21907_ (.A(_19005_),
    .B(_18910_),
    .Y(_19006_));
 sky130_fd_sc_hd__and3_1 _21908_ (.A(_19006_),
    .B(_18988_),
    .C(_19003_),
    .X(_03898_));
 sky130_fd_sc_hd__nand2_1 _21909_ (.A(_19001_),
    .B(_19000_),
    .Y(_19007_));
 sky130_fd_sc_hd__and3_1 _21910_ (.A(_19005_),
    .B(_18988_),
    .C(_19007_),
    .X(_03897_));
 sky130_vsdinv _21911_ (.A(\count_instr[28] ),
    .Y(_19008_));
 sky130_fd_sc_hd__nor2_2 _21912_ (.A(_18886_),
    .B(_18907_),
    .Y(_19009_));
 sky130_fd_sc_hd__nand2_1 _21913_ (.A(_19009_),
    .B(\count_instr[27] ),
    .Y(_19010_));
 sky130_fd_sc_hd__nor2_1 _21914_ (.A(_19008_),
    .B(_19010_),
    .Y(_19011_));
 sky130_fd_sc_hd__and3_1 _21915_ (.A(_19011_),
    .B(\count_instr[30] ),
    .C(\count_instr[29] ),
    .X(_19012_));
 sky130_fd_sc_hd__o211a_1 _21916_ (.A1(\count_instr[31] ),
    .A2(_19012_),
    .B1(_18866_),
    .C1(_19001_),
    .X(_03896_));
 sky130_vsdinv _21917_ (.A(\count_instr[30] ),
    .Y(_19013_));
 sky130_fd_sc_hd__and4_1 _21918_ (.A(_19009_),
    .B(\count_instr[29] ),
    .C(\count_instr[28] ),
    .D(\count_instr[27] ),
    .X(_19014_));
 sky130_vsdinv _21919_ (.A(_19014_),
    .Y(_19015_));
 sky130_fd_sc_hd__a211oi_2 _21920_ (.A1(_19013_),
    .A2(_19015_),
    .B1(_18569_),
    .C1(_19012_),
    .Y(_03895_));
 sky130_fd_sc_hd__o211a_1 _21921_ (.A1(\count_instr[29] ),
    .A2(_19011_),
    .B1(_18866_),
    .C1(_19015_),
    .X(_03894_));
 sky130_fd_sc_hd__or2_1 _21922_ (.A(_18984_),
    .B(_19011_),
    .X(_19016_));
 sky130_fd_sc_hd__a21oi_1 _21923_ (.A1(_19008_),
    .A2(_19010_),
    .B1(_19016_),
    .Y(_03893_));
 sky130_fd_sc_hd__or2_1 _21924_ (.A(\count_instr[27] ),
    .B(_19009_),
    .X(_19017_));
 sky130_fd_sc_hd__and3_1 _21925_ (.A(_19017_),
    .B(_18988_),
    .C(_19010_),
    .X(_03892_));
 sky130_fd_sc_hd__or2_1 _21926_ (.A(_18884_),
    .B(_18907_),
    .X(_19018_));
 sky130_fd_sc_hd__or2_1 _21927_ (.A(_18984_),
    .B(_19009_),
    .X(_19019_));
 sky130_fd_sc_hd__a21oi_1 _21928_ (.A1(_18883_),
    .A2(_19018_),
    .B1(_19019_),
    .Y(_03891_));
 sky130_fd_sc_hd__buf_2 _21929_ (.A(_18331_),
    .X(_19020_));
 sky130_fd_sc_hd__clkbuf_2 _21930_ (.A(_19020_),
    .X(_19021_));
 sky130_fd_sc_hd__nand2_1 _21931_ (.A(_18907_),
    .B(_18884_),
    .Y(_19022_));
 sky130_fd_sc_hd__and3_1 _21932_ (.A(_19018_),
    .B(_19021_),
    .C(_19022_),
    .X(_03890_));
 sky130_fd_sc_hd__nand2_1 _21933_ (.A(_18903_),
    .B(_18906_),
    .Y(_19023_));
 sky130_vsdinv _21934_ (.A(\count_instr[24] ),
    .Y(_19024_));
 sky130_fd_sc_hd__nand2_1 _21935_ (.A(_19023_),
    .B(_19024_),
    .Y(_19025_));
 sky130_fd_sc_hd__and3_1 _21936_ (.A(_19025_),
    .B(_19021_),
    .C(_18907_),
    .X(_03889_));
 sky130_fd_sc_hd__nand2_1 _21937_ (.A(_18903_),
    .B(\count_instr[22] ),
    .Y(_19026_));
 sky130_fd_sc_hd__nand2_1 _21938_ (.A(_19026_),
    .B(_18904_),
    .Y(_19027_));
 sky130_fd_sc_hd__and3_1 _21939_ (.A(_19027_),
    .B(_19021_),
    .C(_19023_),
    .X(_03888_));
 sky130_vsdinv _21940_ (.A(_18903_),
    .Y(_19028_));
 sky130_fd_sc_hd__nand2_1 _21941_ (.A(_19028_),
    .B(_18905_),
    .Y(_19029_));
 sky130_fd_sc_hd__and3_1 _21942_ (.A(_19029_),
    .B(_19021_),
    .C(_19026_),
    .X(_03887_));
 sky130_fd_sc_hd__nand2_1 _21943_ (.A(_18899_),
    .B(\count_instr[19] ),
    .Y(_19030_));
 sky130_fd_sc_hd__nor2_1 _21944_ (.A(_18900_),
    .B(_19030_),
    .Y(_19031_));
 sky130_fd_sc_hd__or2_1 _21945_ (.A(\count_instr[21] ),
    .B(_19031_),
    .X(_19032_));
 sky130_fd_sc_hd__and3_1 _21946_ (.A(_19032_),
    .B(_19021_),
    .C(_19028_),
    .X(_03886_));
 sky130_fd_sc_hd__or2_1 _21947_ (.A(_18984_),
    .B(_19031_),
    .X(_19033_));
 sky130_fd_sc_hd__a21oi_1 _21948_ (.A1(_18900_),
    .A2(_19030_),
    .B1(_19033_),
    .Y(_03885_));
 sky130_vsdinv _21949_ (.A(_18899_),
    .Y(_19034_));
 sky130_fd_sc_hd__nand2_1 _21950_ (.A(_19034_),
    .B(_18901_),
    .Y(_19035_));
 sky130_fd_sc_hd__and3_1 _21951_ (.A(_19035_),
    .B(_19021_),
    .C(_19030_),
    .X(_03884_));
 sky130_vsdinv _21952_ (.A(\count_instr[17] ),
    .Y(_19036_));
 sky130_fd_sc_hd__nand2_1 _21953_ (.A(_18898_),
    .B(\count_instr[16] ),
    .Y(_19037_));
 sky130_fd_sc_hd__nor2_1 _21954_ (.A(_19036_),
    .B(_19037_),
    .Y(_19038_));
 sky130_fd_sc_hd__or2_1 _21955_ (.A(\count_instr[18] ),
    .B(_19038_),
    .X(_19039_));
 sky130_fd_sc_hd__clkbuf_2 _21956_ (.A(_19020_),
    .X(_19040_));
 sky130_fd_sc_hd__and3_1 _21957_ (.A(_19039_),
    .B(_19040_),
    .C(_19034_),
    .X(_03883_));
 sky130_fd_sc_hd__buf_2 _21958_ (.A(_18532_),
    .X(_19041_));
 sky130_fd_sc_hd__or2_1 _21959_ (.A(_19041_),
    .B(_19038_),
    .X(_19042_));
 sky130_fd_sc_hd__a21oi_1 _21960_ (.A1(_19036_),
    .A2(_19037_),
    .B1(_19042_),
    .Y(_03882_));
 sky130_vsdinv _21961_ (.A(_18898_),
    .Y(_19043_));
 sky130_vsdinv _21962_ (.A(\count_instr[16] ),
    .Y(_19044_));
 sky130_fd_sc_hd__nand2_1 _21963_ (.A(_19043_),
    .B(_19044_),
    .Y(_19045_));
 sky130_fd_sc_hd__and3_1 _21964_ (.A(_19045_),
    .B(_19040_),
    .C(_19037_),
    .X(_03881_));
 sky130_fd_sc_hd__a21o_1 _21965_ (.A1(_18897_),
    .A2(\count_instr[14] ),
    .B1(\count_instr[15] ),
    .X(_19046_));
 sky130_fd_sc_hd__and3_1 _21966_ (.A(_19043_),
    .B(_19040_),
    .C(_19046_),
    .X(_03880_));
 sky130_fd_sc_hd__or2_1 _21967_ (.A(\count_instr[14] ),
    .B(_18897_),
    .X(_19047_));
 sky130_fd_sc_hd__nand2_1 _21968_ (.A(_18897_),
    .B(\count_instr[14] ),
    .Y(_19048_));
 sky130_fd_sc_hd__and3_1 _21969_ (.A(_19047_),
    .B(_19040_),
    .C(_19048_),
    .X(_03879_));
 sky130_fd_sc_hd__or2_1 _21970_ (.A(_19041_),
    .B(_18897_),
    .X(_19049_));
 sky130_fd_sc_hd__a21oi_1 _21971_ (.A1(_18890_),
    .A2(_18896_),
    .B1(_19049_),
    .Y(_03878_));
 sky130_vsdinv _21972_ (.A(\count_instr[10] ),
    .Y(_19050_));
 sky130_vsdinv _21973_ (.A(\count_instr[8] ),
    .Y(_19051_));
 sky130_vsdinv _21974_ (.A(\count_instr[7] ),
    .Y(_19052_));
 sky130_vsdinv _21975_ (.A(\count_instr[6] ),
    .Y(_19053_));
 sky130_vsdinv _21976_ (.A(\count_instr[4] ),
    .Y(_19054_));
 sky130_vsdinv _21977_ (.A(\count_instr[0] ),
    .Y(_19055_));
 sky130_vsdinv _21978_ (.A(_18448_),
    .Y(_19056_));
 sky130_fd_sc_hd__nor2_1 _21979_ (.A(_19055_),
    .B(_19056_),
    .Y(_19057_));
 sky130_fd_sc_hd__and3_1 _21980_ (.A(_19057_),
    .B(\count_instr[2] ),
    .C(\count_instr[1] ),
    .X(_19058_));
 sky130_fd_sc_hd__nand2_1 _21981_ (.A(_19058_),
    .B(\count_instr[3] ),
    .Y(_19059_));
 sky130_fd_sc_hd__nor2_1 _21982_ (.A(_19054_),
    .B(_19059_),
    .Y(_19060_));
 sky130_fd_sc_hd__nand2_1 _21983_ (.A(_19060_),
    .B(\count_instr[5] ),
    .Y(_19061_));
 sky130_fd_sc_hd__or3_4 _21984_ (.A(_19052_),
    .B(_19053_),
    .C(_19061_),
    .X(_19062_));
 sky130_fd_sc_hd__nor2_1 _21985_ (.A(_19051_),
    .B(_19062_),
    .Y(_19063_));
 sky130_fd_sc_hd__nand2_1 _21986_ (.A(_19063_),
    .B(\count_instr[9] ),
    .Y(_19064_));
 sky130_fd_sc_hd__or3b_1 _21987_ (.A(_19050_),
    .B(_19064_),
    .C_N(\count_instr[11] ),
    .X(_19065_));
 sky130_vsdinv _21988_ (.A(\count_instr[12] ),
    .Y(_19066_));
 sky130_fd_sc_hd__nand2_1 _21989_ (.A(_19065_),
    .B(_19066_),
    .Y(_19067_));
 sky130_fd_sc_hd__and3_1 _21990_ (.A(_19067_),
    .B(_19040_),
    .C(_18896_),
    .X(_03877_));
 sky130_fd_sc_hd__nor2_1 _21991_ (.A(_19050_),
    .B(_19064_),
    .Y(_19068_));
 sky130_fd_sc_hd__buf_4 _21992_ (.A(_18865_),
    .X(_19069_));
 sky130_fd_sc_hd__o211a_1 _21993_ (.A1(\count_instr[11] ),
    .A2(_19068_),
    .B1(_19069_),
    .C1(_19065_),
    .X(_03876_));
 sky130_fd_sc_hd__or2_1 _21994_ (.A(_19041_),
    .B(_19068_),
    .X(_19070_));
 sky130_fd_sc_hd__a21oi_1 _21995_ (.A1(_19050_),
    .A2(_19064_),
    .B1(_19070_),
    .Y(_03875_));
 sky130_fd_sc_hd__or2_1 _21996_ (.A(\count_instr[9] ),
    .B(_19063_),
    .X(_19071_));
 sky130_fd_sc_hd__and3_1 _21997_ (.A(_19071_),
    .B(_19040_),
    .C(_19064_),
    .X(_03874_));
 sky130_fd_sc_hd__or2_1 _21998_ (.A(_19041_),
    .B(_19063_),
    .X(_19072_));
 sky130_fd_sc_hd__a21oi_1 _21999_ (.A1(_19051_),
    .A2(_19062_),
    .B1(_19072_),
    .Y(_03873_));
 sky130_fd_sc_hd__nor2_1 _22000_ (.A(_19053_),
    .B(_19061_),
    .Y(_19073_));
 sky130_fd_sc_hd__o211a_1 _22001_ (.A1(\count_instr[7] ),
    .A2(_19073_),
    .B1(_19069_),
    .C1(_19062_),
    .X(_03872_));
 sky130_fd_sc_hd__or2_1 _22002_ (.A(_19041_),
    .B(_19073_),
    .X(_19074_));
 sky130_fd_sc_hd__a21oi_1 _22003_ (.A1(_19053_),
    .A2(_19061_),
    .B1(_19074_),
    .Y(_03871_));
 sky130_fd_sc_hd__or2_1 _22004_ (.A(\count_instr[5] ),
    .B(_19060_),
    .X(_19075_));
 sky130_fd_sc_hd__clkbuf_4 _22005_ (.A(_19020_),
    .X(_19076_));
 sky130_fd_sc_hd__and3_1 _22006_ (.A(_19075_),
    .B(_19076_),
    .C(_19061_),
    .X(_03870_));
 sky130_fd_sc_hd__or2_1 _22007_ (.A(_19041_),
    .B(_19060_),
    .X(_19077_));
 sky130_fd_sc_hd__a21oi_1 _22008_ (.A1(_19054_),
    .A2(_19059_),
    .B1(_19077_),
    .Y(_03869_));
 sky130_vsdinv _22009_ (.A(_19058_),
    .Y(_19078_));
 sky130_vsdinv _22010_ (.A(\count_instr[3] ),
    .Y(_19079_));
 sky130_fd_sc_hd__nand2_1 _22011_ (.A(_19078_),
    .B(_19079_),
    .Y(_19080_));
 sky130_fd_sc_hd__and3_1 _22012_ (.A(_19080_),
    .B(_19076_),
    .C(_19059_),
    .X(_03868_));
 sky130_vsdinv _22013_ (.A(\count_instr[1] ),
    .Y(_19081_));
 sky130_vsdinv _22014_ (.A(_19057_),
    .Y(_19082_));
 sky130_fd_sc_hd__nor2_1 _22015_ (.A(_19081_),
    .B(_19082_),
    .Y(_19083_));
 sky130_fd_sc_hd__o211a_1 _22016_ (.A1(\count_instr[2] ),
    .A2(_19083_),
    .B1(_19069_),
    .C1(_19078_),
    .X(_03867_));
 sky130_fd_sc_hd__o21ai_1 _22017_ (.A1(\count_instr[1] ),
    .A2(_19057_),
    .B1(_18935_),
    .Y(_19084_));
 sky130_fd_sc_hd__nor2_1 _22018_ (.A(_19084_),
    .B(_19083_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _22019_ (.A(_19056_),
    .B(_19055_),
    .Y(_19085_));
 sky130_fd_sc_hd__and3_1 _22020_ (.A(_19082_),
    .B(_19076_),
    .C(_19085_),
    .X(_03865_));
 sky130_fd_sc_hd__nor2_1 _22021_ (.A(\cpu_state[1] ),
    .B(net508),
    .Y(_00315_));
 sky130_fd_sc_hd__or3b_4 _22022_ (.A(_00315_),
    .B(_18524_),
    .C_N(_18340_),
    .X(_19086_));
 sky130_vsdinv _22023_ (.A(_19086_),
    .Y(_19087_));
 sky130_fd_sc_hd__clkbuf_2 _22024_ (.A(_19087_),
    .X(_19088_));
 sky130_fd_sc_hd__clkbuf_2 _22025_ (.A(_19088_),
    .X(_19089_));
 sky130_fd_sc_hd__clkbuf_2 _22026_ (.A(_18543_),
    .X(_19090_));
 sky130_fd_sc_hd__clkbuf_4 _22027_ (.A(_19090_),
    .X(_19091_));
 sky130_fd_sc_hd__buf_2 _22028_ (.A(_19086_),
    .X(_19092_));
 sky130_fd_sc_hd__buf_2 _22029_ (.A(_19092_),
    .X(_19093_));
 sky130_fd_sc_hd__a21o_1 _22030_ (.A1(_19091_),
    .A2(_18439_),
    .B1(_19093_),
    .X(_19094_));
 sky130_fd_sc_hd__o211a_1 _22031_ (.A1(net126),
    .A2(_19089_),
    .B1(_19069_),
    .C1(_19094_),
    .X(_03864_));
 sky130_fd_sc_hd__clkbuf_2 _22032_ (.A(_18543_),
    .X(_19095_));
 sky130_fd_sc_hd__buf_2 _22033_ (.A(_19086_),
    .X(_19096_));
 sky130_fd_sc_hd__a31o_1 _22034_ (.A1(_18434_),
    .A2(_19095_),
    .A3(\irq_pending[30] ),
    .B1(_19096_),
    .X(_19097_));
 sky130_fd_sc_hd__o211a_1 _22035_ (.A1(net125),
    .A2(_19089_),
    .B1(_19069_),
    .C1(_19097_),
    .X(_03863_));
 sky130_fd_sc_hd__a21o_1 _22036_ (.A1(_19091_),
    .A2(_18437_),
    .B1(_19093_),
    .X(_19098_));
 sky130_fd_sc_hd__o211a_1 _22037_ (.A1(net123),
    .A2(_19089_),
    .B1(_19069_),
    .C1(_19098_),
    .X(_03862_));
 sky130_fd_sc_hd__buf_2 _22038_ (.A(_18865_),
    .X(_19099_));
 sky130_fd_sc_hd__buf_2 _22039_ (.A(_18543_),
    .X(_19100_));
 sky130_fd_sc_hd__a31o_1 _22040_ (.A1(_18435_),
    .A2(_19100_),
    .A3(\irq_pending[28] ),
    .B1(_19096_),
    .X(_19101_));
 sky130_fd_sc_hd__o211a_1 _22041_ (.A1(net122),
    .A2(_19089_),
    .B1(_19099_),
    .C1(_19101_),
    .X(_03861_));
 sky130_fd_sc_hd__a21o_1 _22042_ (.A1(_19091_),
    .A2(_18403_),
    .B1(_19093_),
    .X(_19102_));
 sky130_fd_sc_hd__o211a_1 _22043_ (.A1(net121),
    .A2(_19089_),
    .B1(_19099_),
    .C1(_19102_),
    .X(_03860_));
 sky130_fd_sc_hd__a21o_1 _22044_ (.A1(_19091_),
    .A2(_18401_),
    .B1(_19093_),
    .X(_19103_));
 sky130_fd_sc_hd__o211a_1 _22045_ (.A1(net120),
    .A2(_19089_),
    .B1(_19099_),
    .C1(_19103_),
    .X(_03859_));
 sky130_fd_sc_hd__buf_2 _22046_ (.A(_19088_),
    .X(_19104_));
 sky130_fd_sc_hd__a31o_1 _22047_ (.A1(_18397_),
    .A2(_19100_),
    .A3(\irq_pending[25] ),
    .B1(_19096_),
    .X(_19105_));
 sky130_fd_sc_hd__o211a_1 _22048_ (.A1(net119),
    .A2(_19104_),
    .B1(_19099_),
    .C1(_19105_),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_4 _22049_ (.A(_18542_),
    .X(_19106_));
 sky130_fd_sc_hd__buf_2 _22050_ (.A(_19106_),
    .X(_19107_));
 sky130_fd_sc_hd__a21o_1 _22051_ (.A1(_19107_),
    .A2(_18399_),
    .B1(_19093_),
    .X(_19108_));
 sky130_fd_sc_hd__o211a_1 _22052_ (.A1(net118),
    .A2(_19104_),
    .B1(_19099_),
    .C1(_19108_),
    .X(_03857_));
 sky130_fd_sc_hd__a21o_1 _22053_ (.A1(_19107_),
    .A2(_18424_),
    .B1(_19093_),
    .X(_19109_));
 sky130_fd_sc_hd__o211a_1 _22054_ (.A1(net117),
    .A2(_19104_),
    .B1(_19099_),
    .C1(_19109_),
    .X(_03856_));
 sky130_fd_sc_hd__buf_2 _22055_ (.A(_18865_),
    .X(_19110_));
 sky130_fd_sc_hd__clkbuf_2 _22056_ (.A(_19092_),
    .X(_19111_));
 sky130_fd_sc_hd__a21o_1 _22057_ (.A1(_19107_),
    .A2(_18422_),
    .B1(_19111_),
    .X(_19112_));
 sky130_fd_sc_hd__o211a_1 _22058_ (.A1(net116),
    .A2(_19104_),
    .B1(_19110_),
    .C1(_19112_),
    .X(_03855_));
 sky130_fd_sc_hd__buf_2 _22059_ (.A(_19092_),
    .X(_19113_));
 sky130_fd_sc_hd__a31o_1 _22060_ (.A1(_18421_),
    .A2(_19100_),
    .A3(\irq_pending[21] ),
    .B1(_19113_),
    .X(_19114_));
 sky130_fd_sc_hd__o211a_1 _22061_ (.A1(net115),
    .A2(_19104_),
    .B1(_19110_),
    .C1(_19114_),
    .X(_03854_));
 sky130_fd_sc_hd__a21o_1 _22062_ (.A1(_19107_),
    .A2(_18426_),
    .B1(_19111_),
    .X(_19115_));
 sky130_fd_sc_hd__o211a_1 _22063_ (.A1(net114),
    .A2(_19104_),
    .B1(_19110_),
    .C1(_19115_),
    .X(_03853_));
 sky130_fd_sc_hd__buf_2 _22064_ (.A(_19088_),
    .X(_19116_));
 sky130_fd_sc_hd__a21o_1 _22065_ (.A1(_19107_),
    .A2(_18391_),
    .B1(_19111_),
    .X(_19117_));
 sky130_fd_sc_hd__o211a_1 _22066_ (.A1(net112),
    .A2(_19116_),
    .B1(_19110_),
    .C1(_19117_),
    .X(_03852_));
 sky130_fd_sc_hd__a21o_1 _22067_ (.A1(_19107_),
    .A2(_18395_),
    .B1(_19111_),
    .X(_19118_));
 sky130_fd_sc_hd__o211a_1 _22068_ (.A1(net111),
    .A2(_19116_),
    .B1(_19110_),
    .C1(_19118_),
    .X(_03851_));
 sky130_fd_sc_hd__a31o_1 _22069_ (.A1(_18390_),
    .A2(_19100_),
    .A3(\irq_pending[17] ),
    .B1(_19113_),
    .X(_19119_));
 sky130_fd_sc_hd__o211a_1 _22070_ (.A1(net110),
    .A2(_19116_),
    .B1(_19110_),
    .C1(_19119_),
    .X(_03850_));
 sky130_fd_sc_hd__buf_2 _22071_ (.A(_18865_),
    .X(_19120_));
 sky130_fd_sc_hd__clkbuf_2 _22072_ (.A(_19106_),
    .X(_19121_));
 sky130_fd_sc_hd__a21o_1 _22073_ (.A1(_19121_),
    .A2(_18393_),
    .B1(_19111_),
    .X(_19122_));
 sky130_fd_sc_hd__o211a_1 _22074_ (.A1(net109),
    .A2(_19116_),
    .B1(_19120_),
    .C1(_19122_),
    .X(_03849_));
 sky130_fd_sc_hd__a21o_1 _22075_ (.A1(_19121_),
    .A2(_18431_),
    .B1(_19111_),
    .X(_19123_));
 sky130_fd_sc_hd__o211a_1 _22076_ (.A1(net108),
    .A2(_19116_),
    .B1(_19120_),
    .C1(_19123_),
    .X(_03848_));
 sky130_fd_sc_hd__a31o_1 _22077_ (.A1(_18428_),
    .A2(_19100_),
    .A3(\irq_pending[14] ),
    .B1(_19113_),
    .X(_19124_));
 sky130_fd_sc_hd__o211a_1 _22078_ (.A1(net107),
    .A2(_19116_),
    .B1(_19120_),
    .C1(_19124_),
    .X(_03847_));
 sky130_fd_sc_hd__clkbuf_2 _22079_ (.A(_19088_),
    .X(_19125_));
 sky130_fd_sc_hd__clkbuf_2 _22080_ (.A(_19092_),
    .X(_19126_));
 sky130_fd_sc_hd__a21o_1 _22081_ (.A1(_19121_),
    .A2(_18430_),
    .B1(_19126_),
    .X(_19127_));
 sky130_fd_sc_hd__o211a_1 _22082_ (.A1(net106),
    .A2(_19125_),
    .B1(_19120_),
    .C1(_19127_),
    .X(_03846_));
 sky130_fd_sc_hd__a31o_1 _22083_ (.A1(_18429_),
    .A2(_19100_),
    .A3(\irq_pending[12] ),
    .B1(_19113_),
    .X(_19128_));
 sky130_fd_sc_hd__o211a_1 _22084_ (.A1(net105),
    .A2(_19125_),
    .B1(_19120_),
    .C1(_19128_),
    .X(_03845_));
 sky130_fd_sc_hd__a21o_1 _22085_ (.A1(_19121_),
    .A2(_18409_),
    .B1(_19126_),
    .X(_19129_));
 sky130_fd_sc_hd__o211a_1 _22086_ (.A1(net104),
    .A2(_19125_),
    .B1(_19120_),
    .C1(_19129_),
    .X(_03844_));
 sky130_fd_sc_hd__clkbuf_2 _22087_ (.A(_18865_),
    .X(_19130_));
 sky130_fd_sc_hd__buf_2 _22088_ (.A(_18543_),
    .X(_19131_));
 sky130_fd_sc_hd__a31o_1 _22089_ (.A1(_18405_),
    .A2(_19131_),
    .A3(\irq_pending[10] ),
    .B1(_19113_),
    .X(_19132_));
 sky130_fd_sc_hd__o211a_1 _22090_ (.A1(net103),
    .A2(_19125_),
    .B1(_19130_),
    .C1(_19132_),
    .X(_03843_));
 sky130_fd_sc_hd__a21o_1 _22091_ (.A1(_19121_),
    .A2(_18407_),
    .B1(_19126_),
    .X(_19133_));
 sky130_fd_sc_hd__o211a_1 _22092_ (.A1(net133),
    .A2(_19125_),
    .B1(_19130_),
    .C1(_19133_),
    .X(_03842_));
 sky130_fd_sc_hd__a31o_1 _22093_ (.A1(_18406_),
    .A2(_19131_),
    .A3(\irq_pending[8] ),
    .B1(_19113_),
    .X(_19134_));
 sky130_fd_sc_hd__o211a_1 _22094_ (.A1(net132),
    .A2(_19125_),
    .B1(_19130_),
    .C1(_19134_),
    .X(_03841_));
 sky130_fd_sc_hd__clkbuf_2 _22095_ (.A(_19087_),
    .X(_19135_));
 sky130_fd_sc_hd__a21o_1 _22096_ (.A1(_19121_),
    .A2(_18388_),
    .B1(_19126_),
    .X(_19136_));
 sky130_fd_sc_hd__o211a_1 _22097_ (.A1(net131),
    .A2(_19135_),
    .B1(_19130_),
    .C1(_19136_),
    .X(_03840_));
 sky130_fd_sc_hd__a31o_1 _22098_ (.A1(_18382_),
    .A2(_19131_),
    .A3(\irq_pending[6] ),
    .B1(_19092_),
    .X(_19137_));
 sky130_fd_sc_hd__o211a_1 _22099_ (.A1(net130),
    .A2(_19135_),
    .B1(_19130_),
    .C1(_19137_),
    .X(_03839_));
 sky130_fd_sc_hd__a21o_1 _22100_ (.A1(_19095_),
    .A2(_18386_),
    .B1(_19126_),
    .X(_19138_));
 sky130_fd_sc_hd__o211a_1 _22101_ (.A1(net129),
    .A2(_19135_),
    .B1(_19130_),
    .C1(_19138_),
    .X(_03838_));
 sky130_fd_sc_hd__buf_4 _22102_ (.A(_18332_),
    .X(_19139_));
 sky130_fd_sc_hd__a21o_1 _22103_ (.A1(_19095_),
    .A2(_18384_),
    .B1(_19126_),
    .X(_19140_));
 sky130_fd_sc_hd__o211a_1 _22104_ (.A1(net128),
    .A2(_19135_),
    .B1(_19139_),
    .C1(_19140_),
    .X(_03837_));
 sky130_fd_sc_hd__a21o_1 _22105_ (.A1(_19095_),
    .A2(_18419_),
    .B1(_19096_),
    .X(_19141_));
 sky130_fd_sc_hd__o211a_1 _22106_ (.A1(net127),
    .A2(_19135_),
    .B1(_19139_),
    .C1(_19141_),
    .X(_03836_));
 sky130_fd_sc_hd__a31o_1 _22107_ (.A1(_18623_),
    .A2(_19131_),
    .A3(\irq_pending[2] ),
    .B1(_19092_),
    .X(_19142_));
 sky130_fd_sc_hd__o211a_1 _22108_ (.A1(net124),
    .A2(_19135_),
    .B1(_19139_),
    .C1(_19142_),
    .X(_03835_));
 sky130_fd_sc_hd__a21o_1 _22109_ (.A1(_19095_),
    .A2(_18417_),
    .B1(_19096_),
    .X(_19143_));
 sky130_fd_sc_hd__o211a_1 _22110_ (.A1(net113),
    .A2(_19088_),
    .B1(_19139_),
    .C1(_19143_),
    .X(_03834_));
 sky130_fd_sc_hd__a21o_1 _22111_ (.A1(_19095_),
    .A2(_18415_),
    .B1(_19096_),
    .X(_19144_));
 sky130_fd_sc_hd__o211a_1 _22112_ (.A1(net102),
    .A2(_19088_),
    .B1(_19139_),
    .C1(_19144_),
    .X(_03833_));
 sky130_fd_sc_hd__nor2_8 _22113_ (.A(instr_ecall_ebreak),
    .B(pcpi_timeout),
    .Y(_00311_));
 sky130_fd_sc_hd__and2_1 _22114_ (.A(_00311_),
    .B(_18462_),
    .X(_19145_));
 sky130_fd_sc_hd__nor2_2 _22115_ (.A(_18520_),
    .B(_18547_),
    .Y(_19146_));
 sky130_vsdinv _22116_ (.A(_19146_),
    .Y(_19147_));
 sky130_fd_sc_hd__or2_1 _22117_ (.A(net370),
    .B(_19146_),
    .X(_19148_));
 sky130_fd_sc_hd__o211a_1 _22118_ (.A1(_19145_),
    .A2(_19147_),
    .B1(_19139_),
    .C1(_19148_),
    .X(_03832_));
 sky130_fd_sc_hd__o21ai_1 _22119_ (.A1(_00290_),
    .A2(_18316_),
    .B1(net237),
    .Y(_19149_));
 sky130_fd_sc_hd__a21o_1 _22120_ (.A1(_18633_),
    .A2(_19149_),
    .B1(net408),
    .X(_19150_));
 sky130_fd_sc_hd__or2b_1 _22121_ (.A(net511),
    .B_N(net237),
    .X(_19151_));
 sky130_fd_sc_hd__a21oi_1 _22122_ (.A1(_19150_),
    .A2(_19151_),
    .B1(_18683_),
    .Y(_03831_));
 sky130_fd_sc_hd__or4_4 _22123_ (.A(\irq_pending[25] ),
    .B(\irq_pending[24] ),
    .C(\irq_pending[27] ),
    .D(\irq_pending[26] ),
    .X(_19152_));
 sky130_fd_sc_hd__or4_4 _22124_ (.A(\irq_pending[21] ),
    .B(\irq_pending[20] ),
    .C(\irq_pending[23] ),
    .D(\irq_pending[22] ),
    .X(_19153_));
 sky130_fd_sc_hd__or4_4 _22125_ (.A(\irq_pending[17] ),
    .B(\irq_pending[16] ),
    .C(\irq_pending[19] ),
    .D(\irq_pending[18] ),
    .X(_19154_));
 sky130_fd_sc_hd__or4_4 _22126_ (.A(\irq_pending[29] ),
    .B(\irq_pending[28] ),
    .C(\irq_pending[31] ),
    .D(\irq_pending[30] ),
    .X(_19155_));
 sky130_fd_sc_hd__or4_4 _22127_ (.A(_19152_),
    .B(_19153_),
    .C(_19154_),
    .D(_19155_),
    .X(_19156_));
 sky130_fd_sc_hd__or4_4 _22128_ (.A(\irq_pending[9] ),
    .B(\irq_pending[8] ),
    .C(\irq_pending[11] ),
    .D(\irq_pending[10] ),
    .X(_19157_));
 sky130_fd_sc_hd__or4_4 _22129_ (.A(\irq_pending[5] ),
    .B(\irq_pending[4] ),
    .C(\irq_pending[7] ),
    .D(\irq_pending[6] ),
    .X(_19158_));
 sky130_fd_sc_hd__or4_4 _22130_ (.A(\irq_pending[1] ),
    .B(\irq_pending[0] ),
    .C(\irq_pending[3] ),
    .D(\irq_pending[2] ),
    .X(_19159_));
 sky130_fd_sc_hd__or4_4 _22131_ (.A(\irq_pending[13] ),
    .B(\irq_pending[12] ),
    .C(\irq_pending[15] ),
    .D(\irq_pending[14] ),
    .X(_19160_));
 sky130_fd_sc_hd__or4_4 _22132_ (.A(_19157_),
    .B(_19158_),
    .C(_19159_),
    .D(_19160_),
    .X(_19161_));
 sky130_fd_sc_hd__nor2_8 _22133_ (.A(_19156_),
    .B(_19161_),
    .Y(_02410_));
 sky130_vsdinv _22134_ (.A(_00309_),
    .Y(_19162_));
 sky130_fd_sc_hd__nor2_1 _22135_ (.A(_18309_),
    .B(_18446_),
    .Y(_19163_));
 sky130_vsdinv _22136_ (.A(_19163_),
    .Y(_19164_));
 sky130_fd_sc_hd__nor2_1 _22137_ (.A(_19162_),
    .B(_19164_),
    .Y(_19165_));
 sky130_fd_sc_hd__and3_1 _22138_ (.A(_19165_),
    .B(_18793_),
    .C(_02410_),
    .X(_03830_));
 sky130_fd_sc_hd__or4_1 _22139_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(instr_sltu),
    .C(instr_slt),
    .D(_18514_),
    .X(_19166_));
 sky130_fd_sc_hd__and3_1 _22140_ (.A(_19166_),
    .B(_19076_),
    .C(_18712_),
    .X(_03829_));
 sky130_fd_sc_hd__nor2_1 _22141_ (.A(mem_do_prefetch),
    .B(_18322_),
    .Y(_19167_));
 sky130_fd_sc_hd__and3_1 _22142_ (.A(_19167_),
    .B(_18330_),
    .C(_18553_),
    .X(_19168_));
 sky130_fd_sc_hd__buf_1 _22143_ (.A(_19168_),
    .X(_03828_));
 sky130_fd_sc_hd__nor2_1 _22144_ (.A(_18534_),
    .B(_18737_),
    .Y(_03827_));
 sky130_fd_sc_hd__and2_1 _22145_ (.A(_18696_),
    .B(_02435_),
    .X(_03826_));
 sky130_fd_sc_hd__and2_1 _22146_ (.A(_18696_),
    .B(_02434_),
    .X(_03825_));
 sky130_fd_sc_hd__and2_1 _22147_ (.A(_18696_),
    .B(_02432_),
    .X(_03824_));
 sky130_fd_sc_hd__buf_1 _22148_ (.A(_18695_),
    .X(_19169_));
 sky130_fd_sc_hd__and2_1 _22149_ (.A(_19169_),
    .B(_02431_),
    .X(_03823_));
 sky130_fd_sc_hd__and2_1 _22150_ (.A(_19169_),
    .B(_02430_),
    .X(_03822_));
 sky130_fd_sc_hd__and2_1 _22151_ (.A(_19169_),
    .B(_02429_),
    .X(_03821_));
 sky130_fd_sc_hd__and2_1 _22152_ (.A(_19169_),
    .B(_02428_),
    .X(_03820_));
 sky130_fd_sc_hd__and2_1 _22153_ (.A(_19169_),
    .B(_02427_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_1 _22154_ (.A(_19169_),
    .B(_02426_),
    .X(_03818_));
 sky130_fd_sc_hd__buf_1 _22155_ (.A(_18695_),
    .X(_19170_));
 sky130_fd_sc_hd__and2_1 _22156_ (.A(_19170_),
    .B(_02425_),
    .X(_03817_));
 sky130_fd_sc_hd__and2_1 _22157_ (.A(_19170_),
    .B(_02424_),
    .X(_03816_));
 sky130_fd_sc_hd__and2_1 _22158_ (.A(_19170_),
    .B(_02423_),
    .X(_03815_));
 sky130_fd_sc_hd__and2_1 _22159_ (.A(_19170_),
    .B(_02421_),
    .X(_03814_));
 sky130_fd_sc_hd__and2_1 _22160_ (.A(_19170_),
    .B(_02420_),
    .X(_03813_));
 sky130_fd_sc_hd__and2_1 _22161_ (.A(_19170_),
    .B(_02419_),
    .X(_03812_));
 sky130_fd_sc_hd__clkbuf_2 _22162_ (.A(_18695_),
    .X(_19171_));
 sky130_fd_sc_hd__and2_1 _22163_ (.A(_19171_),
    .B(_02418_),
    .X(_03811_));
 sky130_fd_sc_hd__and2_1 _22164_ (.A(_19171_),
    .B(_02417_),
    .X(_03810_));
 sky130_fd_sc_hd__and2_1 _22165_ (.A(_19171_),
    .B(_02416_),
    .X(_03809_));
 sky130_fd_sc_hd__and2_1 _22166_ (.A(_19171_),
    .B(_02415_),
    .X(_03808_));
 sky130_fd_sc_hd__and2_1 _22167_ (.A(_19171_),
    .B(_02414_),
    .X(_03807_));
 sky130_fd_sc_hd__and2_1 _22168_ (.A(_19171_),
    .B(_02413_),
    .X(_03806_));
 sky130_fd_sc_hd__clkbuf_2 _22169_ (.A(_18695_),
    .X(_19172_));
 sky130_fd_sc_hd__and2_1 _22170_ (.A(_19172_),
    .B(_02412_),
    .X(_03805_));
 sky130_fd_sc_hd__and2_1 _22171_ (.A(_19172_),
    .B(_02442_),
    .X(_03804_));
 sky130_fd_sc_hd__and2_1 _22172_ (.A(_19172_),
    .B(_02441_),
    .X(_03803_));
 sky130_fd_sc_hd__and2_1 _22173_ (.A(_19172_),
    .B(_02440_),
    .X(_03802_));
 sky130_fd_sc_hd__and2_1 _22174_ (.A(_19172_),
    .B(_02439_),
    .X(_03801_));
 sky130_fd_sc_hd__and2_1 _22175_ (.A(_19172_),
    .B(_02438_),
    .X(_03800_));
 sky130_fd_sc_hd__clkbuf_4 _22176_ (.A(_18934_),
    .X(_19173_));
 sky130_fd_sc_hd__buf_1 _22177_ (.A(_19173_),
    .X(_19174_));
 sky130_fd_sc_hd__and2_1 _22178_ (.A(_19174_),
    .B(_02437_),
    .X(_03799_));
 sky130_fd_sc_hd__and2_1 _22179_ (.A(_19174_),
    .B(_02436_),
    .X(_03798_));
 sky130_fd_sc_hd__and2_1 _22180_ (.A(_19174_),
    .B(_02433_),
    .X(_03797_));
 sky130_fd_sc_hd__and2_1 _22181_ (.A(_19174_),
    .B(_02422_),
    .X(_03796_));
 sky130_fd_sc_hd__and2_1 _22182_ (.A(_19174_),
    .B(_02411_),
    .X(_03795_));
 sky130_vsdinv _22183_ (.A(\count_cycle[63] ),
    .Y(_19175_));
 sky130_fd_sc_hd__nand2_2 _22184_ (.A(\count_cycle[56] ),
    .B(\count_cycle[57] ),
    .Y(_19176_));
 sky130_fd_sc_hd__nand2_1 _22185_ (.A(\count_cycle[58] ),
    .B(\count_cycle[59] ),
    .Y(_19177_));
 sky130_fd_sc_hd__and3_1 _22186_ (.A(\count_cycle[41] ),
    .B(\count_cycle[42] ),
    .C(\count_cycle[43] ),
    .X(_19178_));
 sky130_vsdinv _22187_ (.A(_19178_),
    .Y(_19179_));
 sky130_vsdinv _22188_ (.A(\count_cycle[37] ),
    .Y(_19180_));
 sky130_fd_sc_hd__nand2_2 _22189_ (.A(\count_cycle[35] ),
    .B(\count_cycle[36] ),
    .Y(_19181_));
 sky130_fd_sc_hd__inv_2 _22190_ (.A(\count_cycle[24] ),
    .Y(_01992_));
 sky130_fd_sc_hd__inv_2 _22191_ (.A(\count_cycle[20] ),
    .Y(_01956_));
 sky130_fd_sc_hd__inv_2 _22192_ (.A(\count_cycle[18] ),
    .Y(_01938_));
 sky130_fd_sc_hd__inv_2 _22193_ (.A(\count_cycle[17] ),
    .Y(_01929_));
 sky130_fd_sc_hd__inv_2 _22194_ (.A(\count_cycle[15] ),
    .Y(_01911_));
 sky130_fd_sc_hd__inv_2 _22195_ (.A(\count_cycle[14] ),
    .Y(_01898_));
 sky130_fd_sc_hd__inv_2 _22196_ (.A(\count_cycle[12] ),
    .Y(_01872_));
 sky130_fd_sc_hd__inv_2 _22197_ (.A(\count_cycle[10] ),
    .Y(_01846_));
 sky130_fd_sc_hd__inv_2 _22198_ (.A(\count_cycle[9] ),
    .Y(_01833_));
 sky130_fd_sc_hd__inv_2 _22199_ (.A(\count_cycle[7] ),
    .Y(_01806_));
 sky130_fd_sc_hd__inv_2 _22200_ (.A(\count_cycle[8] ),
    .Y(_01820_));
 sky130_fd_sc_hd__inv_2 _22201_ (.A(\count_cycle[5] ),
    .Y(_01780_));
 sky130_fd_sc_hd__inv_2 _22202_ (.A(\count_cycle[3] ),
    .Y(_01754_));
 sky130_fd_sc_hd__nand2_1 _22203_ (.A(\count_cycle[0] ),
    .B(\count_cycle[1] ),
    .Y(_19182_));
 sky130_fd_sc_hd__inv_2 _22204_ (.A(\count_cycle[2] ),
    .Y(_01741_));
 sky130_fd_sc_hd__or2_1 _22205_ (.A(_19182_),
    .B(_01741_),
    .X(_19183_));
 sky130_fd_sc_hd__nor2_1 _22206_ (.A(_01754_),
    .B(_19183_),
    .Y(_19184_));
 sky130_fd_sc_hd__nand2_1 _22207_ (.A(_19184_),
    .B(\count_cycle[4] ),
    .Y(_19185_));
 sky130_fd_sc_hd__nor2_1 _22208_ (.A(_01780_),
    .B(_19185_),
    .Y(_19186_));
 sky130_fd_sc_hd__nand2_1 _22209_ (.A(_19186_),
    .B(\count_cycle[6] ),
    .Y(_19187_));
 sky130_fd_sc_hd__or3_1 _22210_ (.A(_01806_),
    .B(_01820_),
    .C(_19187_),
    .X(_19188_));
 sky130_fd_sc_hd__or2_1 _22211_ (.A(_01833_),
    .B(_19188_),
    .X(_19189_));
 sky130_fd_sc_hd__nor2_2 _22212_ (.A(_01846_),
    .B(_19189_),
    .Y(_19190_));
 sky130_fd_sc_hd__nand2_4 _22213_ (.A(_19190_),
    .B(\count_cycle[11] ),
    .Y(_19191_));
 sky130_fd_sc_hd__nor2_1 _22214_ (.A(_01872_),
    .B(_19191_),
    .Y(_19192_));
 sky130_fd_sc_hd__nand2_1 _22215_ (.A(_19192_),
    .B(\count_cycle[13] ),
    .Y(_19193_));
 sky130_fd_sc_hd__or2_1 _22216_ (.A(_01898_),
    .B(_19193_),
    .X(_19194_));
 sky130_fd_sc_hd__nor2_1 _22217_ (.A(_01911_),
    .B(_19194_),
    .Y(_19195_));
 sky130_fd_sc_hd__nand2_1 _22218_ (.A(_19195_),
    .B(\count_cycle[16] ),
    .Y(_19196_));
 sky130_fd_sc_hd__or2_1 _22219_ (.A(_01929_),
    .B(_19196_),
    .X(_19197_));
 sky130_fd_sc_hd__nor2_1 _22220_ (.A(_01938_),
    .B(_19197_),
    .Y(_19198_));
 sky130_fd_sc_hd__nand2_1 _22221_ (.A(_19198_),
    .B(\count_cycle[19] ),
    .Y(_19199_));
 sky130_fd_sc_hd__nor2_2 _22222_ (.A(_01956_),
    .B(_19199_),
    .Y(_19200_));
 sky130_fd_sc_hd__and3_1 _22223_ (.A(\count_cycle[21] ),
    .B(\count_cycle[22] ),
    .C(\count_cycle[23] ),
    .X(_19201_));
 sky130_fd_sc_hd__nand2_1 _22224_ (.A(_19200_),
    .B(_19201_),
    .Y(_19202_));
 sky130_fd_sc_hd__nor2_2 _22225_ (.A(_01992_),
    .B(_19202_),
    .Y(_19203_));
 sky130_fd_sc_hd__and3_1 _22226_ (.A(\count_cycle[28] ),
    .B(\count_cycle[29] ),
    .C(\count_cycle[30] ),
    .X(_19204_));
 sky130_fd_sc_hd__and3_1 _22227_ (.A(_19204_),
    .B(\count_cycle[27] ),
    .C(\count_cycle[31] ),
    .X(_19205_));
 sky130_fd_sc_hd__and4_2 _22228_ (.A(_19203_),
    .B(\count_cycle[25] ),
    .C(\count_cycle[26] ),
    .D(_19205_),
    .X(_19206_));
 sky130_vsdinv _22229_ (.A(\count_cycle[33] ),
    .Y(_19207_));
 sky130_vsdinv _22230_ (.A(\count_cycle[34] ),
    .Y(_19208_));
 sky130_fd_sc_hd__nor2_2 _22231_ (.A(_19207_),
    .B(_19208_),
    .Y(_19209_));
 sky130_fd_sc_hd__nand3_4 _22232_ (.A(_19206_),
    .B(\count_cycle[32] ),
    .C(_19209_),
    .Y(_19210_));
 sky130_fd_sc_hd__nor3_4 _22233_ (.A(_19180_),
    .B(_19181_),
    .C(_19210_),
    .Y(_19211_));
 sky130_vsdinv _22234_ (.A(\count_cycle[38] ),
    .Y(_19212_));
 sky130_vsdinv _22235_ (.A(\count_cycle[39] ),
    .Y(_19213_));
 sky130_fd_sc_hd__nor2_2 _22236_ (.A(_19212_),
    .B(_19213_),
    .Y(_19214_));
 sky130_fd_sc_hd__nand3_4 _22237_ (.A(_19211_),
    .B(\count_cycle[40] ),
    .C(_19214_),
    .Y(_19215_));
 sky130_vsdinv _22238_ (.A(\count_cycle[48] ),
    .Y(_19216_));
 sky130_vsdinv _22239_ (.A(\count_cycle[44] ),
    .Y(_19217_));
 sky130_vsdinv _22240_ (.A(\count_cycle[45] ),
    .Y(_19218_));
 sky130_vsdinv _22241_ (.A(\count_cycle[46] ),
    .Y(_19219_));
 sky130_vsdinv _22242_ (.A(\count_cycle[47] ),
    .Y(_19220_));
 sky130_fd_sc_hd__or4_4 _22243_ (.A(_19217_),
    .B(_19218_),
    .C(_19219_),
    .D(_19220_),
    .X(_19221_));
 sky130_fd_sc_hd__nor2_1 _22244_ (.A(_19216_),
    .B(_19221_),
    .Y(_19222_));
 sky130_fd_sc_hd__nor3b_4 _22245_ (.A(_19179_),
    .B(_19215_),
    .C_N(_19222_),
    .Y(_19223_));
 sky130_vsdinv _22246_ (.A(\count_cycle[49] ),
    .Y(_19224_));
 sky130_vsdinv _22247_ (.A(\count_cycle[50] ),
    .Y(_19225_));
 sky130_fd_sc_hd__nor2_4 _22248_ (.A(_19224_),
    .B(_19225_),
    .Y(_19226_));
 sky130_fd_sc_hd__and3_1 _22249_ (.A(\count_cycle[51] ),
    .B(\count_cycle[52] ),
    .C(\count_cycle[53] ),
    .X(_19227_));
 sky130_fd_sc_hd__and3_1 _22250_ (.A(_19227_),
    .B(\count_cycle[54] ),
    .C(\count_cycle[55] ),
    .X(_19228_));
 sky130_fd_sc_hd__nand3_4 _22251_ (.A(_19223_),
    .B(_19226_),
    .C(_19228_),
    .Y(_19229_));
 sky130_fd_sc_hd__nor3_4 _22252_ (.A(_19176_),
    .B(_19177_),
    .C(_19229_),
    .Y(_19230_));
 sky130_fd_sc_hd__clkbuf_2 _22253_ (.A(_19230_),
    .X(_19231_));
 sky130_fd_sc_hd__and2_1 _22254_ (.A(\count_cycle[60] ),
    .B(\count_cycle[61] ),
    .X(_19232_));
 sky130_fd_sc_hd__nand3_1 _22255_ (.A(_19231_),
    .B(\count_cycle[62] ),
    .C(_19232_),
    .Y(_19233_));
 sky130_fd_sc_hd__a41o_1 _22256_ (.A1(_19230_),
    .A2(\count_cycle[62] ),
    .A3(\count_cycle[63] ),
    .A4(_19232_),
    .B1(_18869_),
    .X(_19234_));
 sky130_fd_sc_hd__a21oi_1 _22257_ (.A1(_19175_),
    .A2(_19233_),
    .B1(_19234_),
    .Y(_03794_));
 sky130_fd_sc_hd__a21oi_1 _22258_ (.A1(_19231_),
    .A2(_19232_),
    .B1(\count_cycle[62] ),
    .Y(_19235_));
 sky130_fd_sc_hd__nor3b_1 _22259_ (.A(_18870_),
    .B(_19235_),
    .C_N(_19233_),
    .Y(_03793_));
 sky130_vsdinv _22260_ (.A(\count_cycle[61] ),
    .Y(_19236_));
 sky130_fd_sc_hd__nand2_1 _22261_ (.A(_19231_),
    .B(\count_cycle[60] ),
    .Y(_19237_));
 sky130_fd_sc_hd__a21o_1 _22262_ (.A1(_19231_),
    .A2(_19232_),
    .B1(_18533_),
    .X(_19238_));
 sky130_fd_sc_hd__a21oi_1 _22263_ (.A1(_19236_),
    .A2(_19237_),
    .B1(_19238_),
    .Y(_03792_));
 sky130_fd_sc_hd__nor2_1 _22264_ (.A(\count_cycle[60] ),
    .B(_19231_),
    .Y(_19239_));
 sky130_fd_sc_hd__nor3b_1 _22265_ (.A(_18870_),
    .B(_19239_),
    .C_N(_19237_),
    .Y(_03791_));
 sky130_fd_sc_hd__nor2_1 _22266_ (.A(_19176_),
    .B(_19229_),
    .Y(_19240_));
 sky130_fd_sc_hd__and2_1 _22267_ (.A(_19240_),
    .B(\count_cycle[58] ),
    .X(_19241_));
 sky130_fd_sc_hd__nor2_1 _22268_ (.A(_18598_),
    .B(_19231_),
    .Y(_19242_));
 sky130_fd_sc_hd__o21a_1 _22269_ (.A1(\count_cycle[59] ),
    .A2(_19241_),
    .B1(_19242_),
    .X(_03790_));
 sky130_fd_sc_hd__nor2_1 _22270_ (.A(\count_cycle[58] ),
    .B(_19240_),
    .Y(_19243_));
 sky130_fd_sc_hd__nor3_1 _22271_ (.A(_18870_),
    .B(_19243_),
    .C(_19241_),
    .Y(_03789_));
 sky130_vsdinv _22272_ (.A(\count_cycle[57] ),
    .Y(_19244_));
 sky130_vsdinv _22273_ (.A(\count_cycle[56] ),
    .Y(_19245_));
 sky130_fd_sc_hd__or2_1 _22274_ (.A(_19245_),
    .B(_19229_),
    .X(_19246_));
 sky130_fd_sc_hd__or2_1 _22275_ (.A(_18589_),
    .B(_19240_),
    .X(_19247_));
 sky130_fd_sc_hd__a21oi_1 _22276_ (.A1(_19244_),
    .A2(_19246_),
    .B1(_19247_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _22277_ (.A(_19229_),
    .B(_19245_),
    .Y(_19248_));
 sky130_fd_sc_hd__and3_1 _22278_ (.A(_19246_),
    .B(_19076_),
    .C(_19248_),
    .X(_03787_));
 sky130_fd_sc_hd__nand2_1 _22279_ (.A(_19223_),
    .B(_19226_),
    .Y(_19249_));
 sky130_vsdinv _22280_ (.A(_19249_),
    .Y(_19250_));
 sky130_fd_sc_hd__clkbuf_2 _22281_ (.A(_19250_),
    .X(_19251_));
 sky130_fd_sc_hd__a31o_1 _22282_ (.A1(_19251_),
    .A2(\count_cycle[54] ),
    .A3(_19227_),
    .B1(\count_cycle[55] ),
    .X(_19252_));
 sky130_fd_sc_hd__and3_1 _22283_ (.A(_19252_),
    .B(_19076_),
    .C(_19229_),
    .X(_03786_));
 sky130_fd_sc_hd__a21oi_1 _22284_ (.A1(_19251_),
    .A2(_19227_),
    .B1(\count_cycle[54] ),
    .Y(_19253_));
 sky130_fd_sc_hd__a31o_1 _22285_ (.A1(_19251_),
    .A2(\count_cycle[54] ),
    .A3(_19227_),
    .B1(_18533_),
    .X(_19254_));
 sky130_fd_sc_hd__nor2_1 _22286_ (.A(_19253_),
    .B(_19254_),
    .Y(_03785_));
 sky130_vsdinv _22287_ (.A(_19227_),
    .Y(_19255_));
 sky130_fd_sc_hd__a31o_1 _22288_ (.A1(_19251_),
    .A2(\count_cycle[51] ),
    .A3(\count_cycle[52] ),
    .B1(\count_cycle[53] ),
    .X(_19256_));
 sky130_fd_sc_hd__o211a_1 _22289_ (.A1(_19249_),
    .A2(_19255_),
    .B1(_18938_),
    .C1(_19256_),
    .X(_03784_));
 sky130_vsdinv _22290_ (.A(\count_cycle[52] ),
    .Y(_19257_));
 sky130_fd_sc_hd__nand2_1 _22291_ (.A(_19251_),
    .B(\count_cycle[51] ),
    .Y(_19258_));
 sky130_fd_sc_hd__a31o_1 _22292_ (.A1(_19251_),
    .A2(\count_cycle[51] ),
    .A3(\count_cycle[52] ),
    .B1(_18869_),
    .X(_19259_));
 sky130_fd_sc_hd__a21oi_1 _22293_ (.A1(_19257_),
    .A2(_19258_),
    .B1(_19259_),
    .Y(_03783_));
 sky130_fd_sc_hd__or2_1 _22294_ (.A(\count_cycle[51] ),
    .B(_19250_),
    .X(_19260_));
 sky130_fd_sc_hd__clkbuf_2 _22295_ (.A(_19020_),
    .X(_19261_));
 sky130_fd_sc_hd__and3_1 _22296_ (.A(_19260_),
    .B(_19261_),
    .C(_19258_),
    .X(_03782_));
 sky130_fd_sc_hd__nand2_1 _22297_ (.A(_19223_),
    .B(\count_cycle[49] ),
    .Y(_19262_));
 sky130_fd_sc_hd__nand2_1 _22298_ (.A(_19262_),
    .B(_19225_),
    .Y(_19263_));
 sky130_fd_sc_hd__and3_1 _22299_ (.A(_19263_),
    .B(_19261_),
    .C(_19249_),
    .X(_03781_));
 sky130_vsdinv _22300_ (.A(_19223_),
    .Y(_19264_));
 sky130_fd_sc_hd__nand2_1 _22301_ (.A(_19264_),
    .B(_19224_),
    .Y(_19265_));
 sky130_fd_sc_hd__and3_1 _22302_ (.A(_19265_),
    .B(_19262_),
    .C(_18938_),
    .X(_03780_));
 sky130_fd_sc_hd__nor2_1 _22303_ (.A(_19179_),
    .B(_19215_),
    .Y(_19266_));
 sky130_vsdinv _22304_ (.A(_19266_),
    .Y(_19267_));
 sky130_fd_sc_hd__or2_1 _22305_ (.A(_19221_),
    .B(_19267_),
    .X(_19268_));
 sky130_fd_sc_hd__nand2_1 _22306_ (.A(_19268_),
    .B(_19216_),
    .Y(_19269_));
 sky130_fd_sc_hd__and3_1 _22307_ (.A(_19269_),
    .B(_19261_),
    .C(_19264_),
    .X(_03779_));
 sky130_fd_sc_hd__nand2_1 _22308_ (.A(_19266_),
    .B(\count_cycle[44] ),
    .Y(_19270_));
 sky130_fd_sc_hd__or3_1 _22309_ (.A(_19218_),
    .B(_19219_),
    .C(_19270_),
    .X(_19271_));
 sky130_fd_sc_hd__nand2_1 _22310_ (.A(_19271_),
    .B(_19220_),
    .Y(_19272_));
 sky130_fd_sc_hd__and3_1 _22311_ (.A(_19272_),
    .B(_19261_),
    .C(_19268_),
    .X(_03778_));
 sky130_fd_sc_hd__or2_1 _22312_ (.A(_19218_),
    .B(_19270_),
    .X(_19273_));
 sky130_fd_sc_hd__nand2_1 _22313_ (.A(_19273_),
    .B(_19219_),
    .Y(_19274_));
 sky130_fd_sc_hd__and3_1 _22314_ (.A(_19274_),
    .B(_19271_),
    .C(_18938_),
    .X(_03777_));
 sky130_fd_sc_hd__nand2_1 _22315_ (.A(_19270_),
    .B(_19218_),
    .Y(_19275_));
 sky130_fd_sc_hd__and3_1 _22316_ (.A(_19273_),
    .B(_19261_),
    .C(_19275_),
    .X(_03776_));
 sky130_fd_sc_hd__nand2_1 _22317_ (.A(_19267_),
    .B(_19217_),
    .Y(_19276_));
 sky130_fd_sc_hd__and3_1 _22318_ (.A(_19276_),
    .B(_19261_),
    .C(_19270_),
    .X(_03775_));
 sky130_vsdinv _22319_ (.A(\count_cycle[42] ),
    .Y(_19277_));
 sky130_vsdinv _22320_ (.A(_19215_),
    .Y(_19278_));
 sky130_fd_sc_hd__nand2_1 _22321_ (.A(_19278_),
    .B(\count_cycle[41] ),
    .Y(_19279_));
 sky130_fd_sc_hd__or2_1 _22322_ (.A(_19277_),
    .B(_19279_),
    .X(_19280_));
 sky130_vsdinv _22323_ (.A(\count_cycle[43] ),
    .Y(_19281_));
 sky130_fd_sc_hd__nand2_1 _22324_ (.A(_19280_),
    .B(_19281_),
    .Y(_19282_));
 sky130_fd_sc_hd__buf_1 _22325_ (.A(_19020_),
    .X(_19283_));
 sky130_fd_sc_hd__and3_1 _22326_ (.A(_19282_),
    .B(_19283_),
    .C(_19267_),
    .X(_03774_));
 sky130_fd_sc_hd__nand2_1 _22327_ (.A(_19279_),
    .B(_19277_),
    .Y(_19284_));
 sky130_fd_sc_hd__and3_1 _22328_ (.A(_19280_),
    .B(_19283_),
    .C(_19284_),
    .X(_03773_));
 sky130_fd_sc_hd__or2_1 _22329_ (.A(\count_cycle[41] ),
    .B(_19278_),
    .X(_19285_));
 sky130_fd_sc_hd__and3_1 _22330_ (.A(_19285_),
    .B(_19283_),
    .C(_19279_),
    .X(_03772_));
 sky130_fd_sc_hd__nand2_1 _22331_ (.A(_19211_),
    .B(_19214_),
    .Y(_19286_));
 sky130_vsdinv _22332_ (.A(\count_cycle[40] ),
    .Y(_19287_));
 sky130_fd_sc_hd__nand2_1 _22333_ (.A(_19286_),
    .B(_19287_),
    .Y(_19288_));
 sky130_fd_sc_hd__and3_1 _22334_ (.A(_19288_),
    .B(_19283_),
    .C(_19215_),
    .X(_03771_));
 sky130_fd_sc_hd__nand2_1 _22335_ (.A(_19211_),
    .B(\count_cycle[38] ),
    .Y(_19289_));
 sky130_fd_sc_hd__nand2_1 _22336_ (.A(_19289_),
    .B(_19213_),
    .Y(_19290_));
 sky130_fd_sc_hd__and3_1 _22337_ (.A(_19290_),
    .B(_19283_),
    .C(_19286_),
    .X(_03770_));
 sky130_vsdinv _22338_ (.A(_19211_),
    .Y(_19291_));
 sky130_fd_sc_hd__nand2_1 _22339_ (.A(_19291_),
    .B(_19212_),
    .Y(_19292_));
 sky130_fd_sc_hd__and3_1 _22340_ (.A(_19292_),
    .B(_19283_),
    .C(_19289_),
    .X(_03769_));
 sky130_fd_sc_hd__nor2_1 _22341_ (.A(_19181_),
    .B(_19210_),
    .Y(_19293_));
 sky130_vsdinv _22342_ (.A(_19293_),
    .Y(_19294_));
 sky130_fd_sc_hd__nand2_1 _22343_ (.A(_19294_),
    .B(_19180_),
    .Y(_19295_));
 sky130_fd_sc_hd__clkbuf_2 _22344_ (.A(_19020_),
    .X(_19296_));
 sky130_fd_sc_hd__and3_1 _22345_ (.A(_19295_),
    .B(_19296_),
    .C(_19291_),
    .X(_03768_));
 sky130_vsdinv _22346_ (.A(\count_cycle[35] ),
    .Y(_19297_));
 sky130_fd_sc_hd__nor2_1 _22347_ (.A(_19297_),
    .B(_19210_),
    .Y(_19298_));
 sky130_vsdinv _22348_ (.A(_19298_),
    .Y(_19299_));
 sky130_vsdinv _22349_ (.A(\count_cycle[36] ),
    .Y(_19300_));
 sky130_fd_sc_hd__nand2_1 _22350_ (.A(_19299_),
    .B(_19300_),
    .Y(_19301_));
 sky130_fd_sc_hd__and3_1 _22351_ (.A(_19301_),
    .B(_19296_),
    .C(_19294_),
    .X(_03767_));
 sky130_fd_sc_hd__nand2_1 _22352_ (.A(_19210_),
    .B(_19297_),
    .Y(_19302_));
 sky130_fd_sc_hd__and3_1 _22353_ (.A(_19299_),
    .B(_19296_),
    .C(_19302_),
    .X(_03766_));
 sky130_vsdinv _22354_ (.A(\count_cycle[32] ),
    .Y(_19303_));
 sky130_vsdinv _22355_ (.A(_19206_),
    .Y(_19304_));
 sky130_fd_sc_hd__nor2_1 _22356_ (.A(_19303_),
    .B(_19304_),
    .Y(_19305_));
 sky130_fd_sc_hd__nand2_1 _22357_ (.A(_19305_),
    .B(\count_cycle[33] ),
    .Y(_19306_));
 sky130_fd_sc_hd__nand2_1 _22358_ (.A(_19306_),
    .B(_19208_),
    .Y(_19307_));
 sky130_fd_sc_hd__and3_1 _22359_ (.A(_19307_),
    .B(_19296_),
    .C(_19210_),
    .X(_03765_));
 sky130_vsdinv _22360_ (.A(_19305_),
    .Y(_19308_));
 sky130_fd_sc_hd__nand2_1 _22361_ (.A(_19308_),
    .B(_19207_),
    .Y(_19309_));
 sky130_fd_sc_hd__and3_1 _22362_ (.A(_19309_),
    .B(_19296_),
    .C(_19306_),
    .X(_03764_));
 sky130_fd_sc_hd__nand2_1 _22363_ (.A(_19304_),
    .B(_19303_),
    .Y(_19310_));
 sky130_fd_sc_hd__and3_1 _22364_ (.A(_19308_),
    .B(_19296_),
    .C(_19310_),
    .X(_03763_));
 sky130_fd_sc_hd__inv_2 _22365_ (.A(\count_cycle[30] ),
    .Y(_02046_));
 sky130_fd_sc_hd__inv_2 _22366_ (.A(\count_cycle[29] ),
    .Y(_02037_));
 sky130_fd_sc_hd__inv_2 _22367_ (.A(\count_cycle[28] ),
    .Y(_02028_));
 sky130_fd_sc_hd__inv_2 _22368_ (.A(\count_cycle[26] ),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _22369_ (.A(_19203_),
    .B(\count_cycle[25] ),
    .Y(_19311_));
 sky130_fd_sc_hd__nor2_1 _22370_ (.A(_02010_),
    .B(_19311_),
    .Y(_19312_));
 sky130_fd_sc_hd__nand2_1 _22371_ (.A(_19312_),
    .B(\count_cycle[27] ),
    .Y(_19313_));
 sky130_fd_sc_hd__or2_1 _22372_ (.A(_02028_),
    .B(_19313_),
    .X(_19314_));
 sky130_fd_sc_hd__or2_1 _22373_ (.A(_02037_),
    .B(_19314_),
    .X(_19315_));
 sky130_fd_sc_hd__or2_1 _22374_ (.A(_02046_),
    .B(_19315_),
    .X(_19316_));
 sky130_fd_sc_hd__inv_2 _22375_ (.A(\count_cycle[31] ),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _22376_ (.A(_19316_),
    .B(_02055_),
    .Y(_19317_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _22377_ (.A(_18934_),
    .X(_19318_));
 sky130_fd_sc_hd__and3_1 _22378_ (.A(_19317_),
    .B(_19318_),
    .C(_19304_),
    .X(_03762_));
 sky130_fd_sc_hd__nand2_1 _22379_ (.A(_19315_),
    .B(_02046_),
    .Y(_19319_));
 sky130_fd_sc_hd__and3_1 _22380_ (.A(_19316_),
    .B(_19318_),
    .C(_19319_),
    .X(_03761_));
 sky130_fd_sc_hd__nand2_1 _22381_ (.A(_19314_),
    .B(_02037_),
    .Y(_19320_));
 sky130_fd_sc_hd__and3_1 _22382_ (.A(_19315_),
    .B(_19318_),
    .C(_19320_),
    .X(_03760_));
 sky130_fd_sc_hd__nand2_1 _22383_ (.A(_19313_),
    .B(_02028_),
    .Y(_19321_));
 sky130_fd_sc_hd__and3_1 _22384_ (.A(_19314_),
    .B(_19318_),
    .C(_19321_),
    .X(_03759_));
 sky130_fd_sc_hd__or2_1 _22385_ (.A(\count_cycle[27] ),
    .B(_19312_),
    .X(_19322_));
 sky130_fd_sc_hd__and3_1 _22386_ (.A(_19322_),
    .B(_19318_),
    .C(_19313_),
    .X(_03758_));
 sky130_fd_sc_hd__or2_1 _22387_ (.A(_18589_),
    .B(_19312_),
    .X(_19323_));
 sky130_fd_sc_hd__a21oi_1 _22388_ (.A1(_02010_),
    .A2(_19311_),
    .B1(_19323_),
    .Y(_03757_));
 sky130_vsdinv _22389_ (.A(_19203_),
    .Y(_19324_));
 sky130_fd_sc_hd__inv_2 _22390_ (.A(\count_cycle[25] ),
    .Y(_02001_));
 sky130_fd_sc_hd__nand2_1 _22391_ (.A(_19324_),
    .B(_02001_),
    .Y(_19325_));
 sky130_fd_sc_hd__and3_1 _22392_ (.A(_19325_),
    .B(_19318_),
    .C(_19311_),
    .X(_03756_));
 sky130_fd_sc_hd__buf_1 _22393_ (.A(_18934_),
    .X(_19326_));
 sky130_fd_sc_hd__nand2_1 _22394_ (.A(_19202_),
    .B(_01992_),
    .Y(_19327_));
 sky130_fd_sc_hd__and3_1 _22395_ (.A(_19324_),
    .B(_19326_),
    .C(_19327_),
    .X(_03755_));
 sky130_fd_sc_hd__inv_2 _22396_ (.A(\count_cycle[22] ),
    .Y(_01974_));
 sky130_fd_sc_hd__nand2_1 _22397_ (.A(_19200_),
    .B(\count_cycle[21] ),
    .Y(_19328_));
 sky130_fd_sc_hd__or2_1 _22398_ (.A(_01974_),
    .B(_19328_),
    .X(_19329_));
 sky130_fd_sc_hd__inv_2 _22399_ (.A(\count_cycle[23] ),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _22400_ (.A(_19329_),
    .B(_01983_),
    .Y(_19330_));
 sky130_fd_sc_hd__and3_1 _22401_ (.A(_19330_),
    .B(_19326_),
    .C(_19202_),
    .X(_03754_));
 sky130_fd_sc_hd__nand2_1 _22402_ (.A(_19328_),
    .B(_01974_),
    .Y(_19331_));
 sky130_fd_sc_hd__and3_1 _22403_ (.A(_19329_),
    .B(_19326_),
    .C(_19331_),
    .X(_03753_));
 sky130_vsdinv _22404_ (.A(_19200_),
    .Y(_19332_));
 sky130_fd_sc_hd__inv_2 _22405_ (.A(\count_cycle[21] ),
    .Y(_01965_));
 sky130_fd_sc_hd__nand2_1 _22406_ (.A(_19332_),
    .B(_01965_),
    .Y(_19333_));
 sky130_fd_sc_hd__and3_1 _22407_ (.A(_19333_),
    .B(_19326_),
    .C(_19328_),
    .X(_03752_));
 sky130_fd_sc_hd__nand2_1 _22408_ (.A(_19199_),
    .B(_01956_),
    .Y(_19334_));
 sky130_fd_sc_hd__and3_1 _22409_ (.A(_19332_),
    .B(_19326_),
    .C(_19334_),
    .X(_03751_));
 sky130_fd_sc_hd__or2_1 _22410_ (.A(\count_cycle[19] ),
    .B(_19198_),
    .X(_19335_));
 sky130_fd_sc_hd__and3_1 _22411_ (.A(_19335_),
    .B(_19326_),
    .C(_19199_),
    .X(_03750_));
 sky130_fd_sc_hd__or2_1 _22412_ (.A(_18589_),
    .B(_19198_),
    .X(_19336_));
 sky130_fd_sc_hd__a21oi_1 _22413_ (.A1(_01938_),
    .A2(_19197_),
    .B1(_19336_),
    .Y(_03749_));
 sky130_fd_sc_hd__clkbuf_2 _22414_ (.A(_18934_),
    .X(_19337_));
 sky130_fd_sc_hd__nand2_1 _22415_ (.A(_19196_),
    .B(_01929_),
    .Y(_19338_));
 sky130_fd_sc_hd__and3_1 _22416_ (.A(_19197_),
    .B(_19337_),
    .C(_19338_),
    .X(_03748_));
 sky130_vsdinv _22417_ (.A(_19195_),
    .Y(_19339_));
 sky130_fd_sc_hd__inv_2 _22418_ (.A(\count_cycle[16] ),
    .Y(_01920_));
 sky130_fd_sc_hd__nand2_1 _22419_ (.A(_19339_),
    .B(_01920_),
    .Y(_19340_));
 sky130_fd_sc_hd__and3_1 _22420_ (.A(_19340_),
    .B(_19337_),
    .C(_19196_),
    .X(_03747_));
 sky130_fd_sc_hd__nand2_1 _22421_ (.A(_19194_),
    .B(_01911_),
    .Y(_19341_));
 sky130_fd_sc_hd__and3_1 _22422_ (.A(_19339_),
    .B(_19337_),
    .C(_19341_),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_1 _22423_ (.A(_19193_),
    .B(_01898_),
    .Y(_19342_));
 sky130_fd_sc_hd__and3_1 _22424_ (.A(_19194_),
    .B(_19337_),
    .C(_19342_),
    .X(_03745_));
 sky130_vsdinv _22425_ (.A(_19192_),
    .Y(_19343_));
 sky130_fd_sc_hd__inv_2 _22426_ (.A(\count_cycle[13] ),
    .Y(_01885_));
 sky130_fd_sc_hd__nand2_1 _22427_ (.A(_19343_),
    .B(_01885_),
    .Y(_19344_));
 sky130_fd_sc_hd__and3_1 _22428_ (.A(_19344_),
    .B(_19337_),
    .C(_19193_),
    .X(_03744_));
 sky130_fd_sc_hd__nand2_1 _22429_ (.A(_19191_),
    .B(_01872_),
    .Y(_19345_));
 sky130_fd_sc_hd__and3_1 _22430_ (.A(_19343_),
    .B(_19337_),
    .C(_19345_),
    .X(_03743_));
 sky130_vsdinv _22431_ (.A(_19190_),
    .Y(_19346_));
 sky130_fd_sc_hd__inv_2 _22432_ (.A(\count_cycle[11] ),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_1 _22433_ (.A(_19346_),
    .B(_01859_),
    .Y(_19347_));
 sky130_fd_sc_hd__clkbuf_2 _22434_ (.A(_18934_),
    .X(_19348_));
 sky130_fd_sc_hd__and3_1 _22435_ (.A(_19347_),
    .B(_19348_),
    .C(_19191_),
    .X(_03742_));
 sky130_fd_sc_hd__nand2_1 _22436_ (.A(_19189_),
    .B(_01846_),
    .Y(_19349_));
 sky130_fd_sc_hd__and3_1 _22437_ (.A(_19346_),
    .B(_19348_),
    .C(_19349_),
    .X(_03741_));
 sky130_fd_sc_hd__nand2_1 _22438_ (.A(_19188_),
    .B(_01833_),
    .Y(_19350_));
 sky130_fd_sc_hd__and3_1 _22439_ (.A(_19189_),
    .B(_19348_),
    .C(_19350_),
    .X(_03740_));
 sky130_fd_sc_hd__or2_1 _22440_ (.A(_01806_),
    .B(_19187_),
    .X(_19351_));
 sky130_fd_sc_hd__nand2_1 _22441_ (.A(_19351_),
    .B(_01820_),
    .Y(_19352_));
 sky130_fd_sc_hd__and3_1 _22442_ (.A(_19352_),
    .B(_19188_),
    .C(_18938_),
    .X(_03739_));
 sky130_fd_sc_hd__nand2_1 _22443_ (.A(_19187_),
    .B(_01806_),
    .Y(_19353_));
 sky130_fd_sc_hd__and3_1 _22444_ (.A(_19351_),
    .B(_19348_),
    .C(_19353_),
    .X(_03738_));
 sky130_vsdinv _22445_ (.A(_19186_),
    .Y(_19354_));
 sky130_fd_sc_hd__inv_2 _22446_ (.A(\count_cycle[6] ),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _22447_ (.A(_19354_),
    .B(_01793_),
    .Y(_19355_));
 sky130_fd_sc_hd__and3_1 _22448_ (.A(_19355_),
    .B(_19348_),
    .C(_19187_),
    .X(_03737_));
 sky130_fd_sc_hd__nand2_1 _22449_ (.A(_19185_),
    .B(_01780_),
    .Y(_19356_));
 sky130_fd_sc_hd__and3_1 _22450_ (.A(_19354_),
    .B(_19348_),
    .C(_19356_),
    .X(_03736_));
 sky130_vsdinv _22451_ (.A(_19184_),
    .Y(_19357_));
 sky130_fd_sc_hd__inv_2 _22452_ (.A(\count_cycle[4] ),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _22453_ (.A(_19357_),
    .B(_01767_),
    .Y(_19358_));
 sky130_fd_sc_hd__and3_1 _22454_ (.A(_19358_),
    .B(_18935_),
    .C(_19185_),
    .X(_03735_));
 sky130_fd_sc_hd__nand2_1 _22455_ (.A(_19183_),
    .B(_01754_),
    .Y(_19359_));
 sky130_fd_sc_hd__and3_1 _22456_ (.A(_19357_),
    .B(_18935_),
    .C(_19359_),
    .X(_03734_));
 sky130_fd_sc_hd__nand2_1 _22457_ (.A(_01741_),
    .B(_19182_),
    .Y(_19360_));
 sky130_fd_sc_hd__and3_1 _22458_ (.A(_19183_),
    .B(_18935_),
    .C(_19360_),
    .X(_03733_));
 sky130_fd_sc_hd__inv_2 _22459_ (.A(\count_cycle[0] ),
    .Y(_02559_));
 sky130_fd_sc_hd__inv_2 _22460_ (.A(\count_cycle[1] ),
    .Y(_01728_));
 sky130_fd_sc_hd__nand2_1 _22461_ (.A(_02559_),
    .B(_01728_),
    .Y(_19361_));
 sky130_fd_sc_hd__and3_1 _22462_ (.A(_19361_),
    .B(_18935_),
    .C(_19182_),
    .X(_03732_));
 sky130_fd_sc_hd__nor2_1 _22463_ (.A(\count_cycle[0] ),
    .B(_18644_),
    .Y(_03731_));
 sky130_vsdinv _22464_ (.A(\cpu_state[0] ),
    .Y(_19362_));
 sky130_fd_sc_hd__nor2_1 _22465_ (.A(_18534_),
    .B(_19362_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor2_1 _22466_ (.A(_18534_),
    .B(_18461_),
    .Y(_03729_));
 sky130_fd_sc_hd__buf_1 _22467_ (.A(\cpuregs_wrdata[31] ),
    .X(_19363_));
 sky130_vsdinv _22468_ (.A(\latched_rd[1] ),
    .Y(_19364_));
 sky130_vsdinv _22469_ (.A(\latched_rd[0] ),
    .Y(_19365_));
 sky130_fd_sc_hd__nand2_2 _22470_ (.A(_19365_),
    .B(_19364_),
    .Y(_19366_));
 sky130_fd_sc_hd__nor2_1 _22471_ (.A(\latched_rd[4] ),
    .B(\latched_rd[2] ),
    .Y(_19367_));
 sky130_vsdinv _22472_ (.A(\latched_rd[3] ),
    .Y(_19368_));
 sky130_fd_sc_hd__nand2_2 _22473_ (.A(_19367_),
    .B(_19368_),
    .Y(_19369_));
 sky130_fd_sc_hd__nor2_8 _22474_ (.A(_18308_),
    .B(_18500_),
    .Y(_19370_));
 sky130_fd_sc_hd__o31a_4 _22475_ (.A1(latched_branch),
    .A2(latched_store),
    .A3(_18536_),
    .B1(_19370_),
    .X(_19371_));
 sky130_fd_sc_hd__o21ai_4 _22476_ (.A1(_19366_),
    .A2(_19369_),
    .B1(_19371_),
    .Y(_19372_));
 sky130_fd_sc_hd__or2_2 _22477_ (.A(_19364_),
    .B(_19372_),
    .X(_19373_));
 sky130_fd_sc_hd__nor2_4 _22478_ (.A(\latched_rd[0] ),
    .B(_19373_),
    .Y(_19374_));
 sky130_vsdinv _22479_ (.A(\latched_rd[4] ),
    .Y(_19375_));
 sky130_fd_sc_hd__and3_1 _22480_ (.A(_19375_),
    .B(_19368_),
    .C(\latched_rd[2] ),
    .X(_19376_));
 sky130_fd_sc_hd__nand2_1 _22481_ (.A(_19374_),
    .B(_19376_),
    .Y(_19377_));
 sky130_fd_sc_hd__clkbuf_8 _22482_ (.A(_19377_),
    .X(_19378_));
 sky130_fd_sc_hd__buf_4 _22483_ (.A(_19378_),
    .X(_19379_));
 sky130_fd_sc_hd__mux2_1 _22484_ (.A0(_19363_),
    .A1(\cpuregs[6][31] ),
    .S(_19379_),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_2 _22485_ (.A(\cpuregs_wrdata[30] ),
    .X(_19380_));
 sky130_fd_sc_hd__mux2_1 _22486_ (.A0(_19380_),
    .A1(\cpuregs[6][30] ),
    .S(_19379_),
    .X(_03726_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _22487_ (.A(\cpuregs_wrdata[29] ),
    .X(_19381_));
 sky130_fd_sc_hd__mux2_1 _22488_ (.A0(_19381_),
    .A1(\cpuregs[6][29] ),
    .S(_19379_),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_2 _22489_ (.A(\cpuregs_wrdata[28] ),
    .X(_19382_));
 sky130_fd_sc_hd__mux2_1 _22490_ (.A0(_19382_),
    .A1(\cpuregs[6][28] ),
    .S(_19379_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_2 _22491_ (.A(\cpuregs_wrdata[27] ),
    .X(_19383_));
 sky130_fd_sc_hd__mux2_1 _22492_ (.A0(_19383_),
    .A1(\cpuregs[6][27] ),
    .S(_19379_),
    .X(_03723_));
 sky130_fd_sc_hd__buf_1 _22493_ (.A(\cpuregs_wrdata[26] ),
    .X(_19384_));
 sky130_fd_sc_hd__mux2_1 _22494_ (.A0(_19384_),
    .A1(\cpuregs[6][26] ),
    .S(_19379_),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_2 _22495_ (.A(\cpuregs_wrdata[25] ),
    .X(_19385_));
 sky130_fd_sc_hd__buf_2 _22496_ (.A(_19378_),
    .X(_19386_));
 sky130_fd_sc_hd__mux2_1 _22497_ (.A0(_19385_),
    .A1(\cpuregs[6][25] ),
    .S(_19386_),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_2 _22498_ (.A(\cpuregs_wrdata[24] ),
    .X(_19387_));
 sky130_fd_sc_hd__mux2_1 _22499_ (.A0(_19387_),
    .A1(\cpuregs[6][24] ),
    .S(_19386_),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_2 _22500_ (.A(\cpuregs_wrdata[23] ),
    .X(_19388_));
 sky130_fd_sc_hd__mux2_1 _22501_ (.A0(_19388_),
    .A1(\cpuregs[6][23] ),
    .S(_19386_),
    .X(_03719_));
 sky130_fd_sc_hd__clkbuf_2 _22502_ (.A(\cpuregs_wrdata[22] ),
    .X(_19389_));
 sky130_fd_sc_hd__mux2_1 _22503_ (.A0(_19389_),
    .A1(\cpuregs[6][22] ),
    .S(_19386_),
    .X(_03718_));
 sky130_fd_sc_hd__clkbuf_2 _22504_ (.A(\cpuregs_wrdata[21] ),
    .X(_19390_));
 sky130_fd_sc_hd__mux2_1 _22505_ (.A0(_19390_),
    .A1(\cpuregs[6][21] ),
    .S(_19386_),
    .X(_03717_));
 sky130_fd_sc_hd__clkbuf_2 _22506_ (.A(\cpuregs_wrdata[20] ),
    .X(_19391_));
 sky130_fd_sc_hd__mux2_1 _22507_ (.A0(_19391_),
    .A1(\cpuregs[6][20] ),
    .S(_19386_),
    .X(_03716_));
 sky130_fd_sc_hd__clkbuf_2 _22508_ (.A(\cpuregs_wrdata[19] ),
    .X(_19392_));
 sky130_fd_sc_hd__clkbuf_4 _22509_ (.A(_19378_),
    .X(_19393_));
 sky130_fd_sc_hd__mux2_1 _22510_ (.A0(_19392_),
    .A1(\cpuregs[6][19] ),
    .S(_19393_),
    .X(_03715_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _22511_ (.A(\cpuregs_wrdata[18] ),
    .X(_19394_));
 sky130_fd_sc_hd__mux2_1 _22512_ (.A0(_19394_),
    .A1(\cpuregs[6][18] ),
    .S(_19393_),
    .X(_03714_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _22513_ (.A(\cpuregs_wrdata[17] ),
    .X(_19395_));
 sky130_fd_sc_hd__mux2_1 _22514_ (.A0(_19395_),
    .A1(\cpuregs[6][17] ),
    .S(_19393_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_2 _22515_ (.A(\cpuregs_wrdata[16] ),
    .X(_19396_));
 sky130_fd_sc_hd__mux2_1 _22516_ (.A0(_19396_),
    .A1(\cpuregs[6][16] ),
    .S(_19393_),
    .X(_03712_));
 sky130_fd_sc_hd__clkbuf_2 _22517_ (.A(\cpuregs_wrdata[15] ),
    .X(_19397_));
 sky130_fd_sc_hd__mux2_1 _22518_ (.A0(_19397_),
    .A1(\cpuregs[6][15] ),
    .S(_19393_),
    .X(_03711_));
 sky130_fd_sc_hd__clkbuf_2 _22519_ (.A(\cpuregs_wrdata[14] ),
    .X(_19398_));
 sky130_fd_sc_hd__mux2_1 _22520_ (.A0(_19398_),
    .A1(\cpuregs[6][14] ),
    .S(_19393_),
    .X(_03710_));
 sky130_fd_sc_hd__clkbuf_2 _22521_ (.A(\cpuregs_wrdata[13] ),
    .X(_19399_));
 sky130_fd_sc_hd__clkbuf_4 _22522_ (.A(_19378_),
    .X(_19400_));
 sky130_fd_sc_hd__mux2_1 _22523_ (.A0(_19399_),
    .A1(\cpuregs[6][13] ),
    .S(_19400_),
    .X(_03709_));
 sky130_fd_sc_hd__clkbuf_2 _22524_ (.A(\cpuregs_wrdata[12] ),
    .X(_19401_));
 sky130_fd_sc_hd__mux2_1 _22525_ (.A0(_19401_),
    .A1(\cpuregs[6][12] ),
    .S(_19400_),
    .X(_03708_));
 sky130_fd_sc_hd__clkbuf_2 _22526_ (.A(\cpuregs_wrdata[11] ),
    .X(_19402_));
 sky130_fd_sc_hd__mux2_1 _22527_ (.A0(_19402_),
    .A1(\cpuregs[6][11] ),
    .S(_19400_),
    .X(_03707_));
 sky130_fd_sc_hd__clkbuf_2 _22528_ (.A(\cpuregs_wrdata[10] ),
    .X(_19403_));
 sky130_fd_sc_hd__mux2_1 _22529_ (.A0(_19403_),
    .A1(\cpuregs[6][10] ),
    .S(_19400_),
    .X(_03706_));
 sky130_fd_sc_hd__clkbuf_2 _22530_ (.A(\cpuregs_wrdata[9] ),
    .X(_19404_));
 sky130_fd_sc_hd__mux2_1 _22531_ (.A0(_19404_),
    .A1(\cpuregs[6][9] ),
    .S(_19400_),
    .X(_03705_));
 sky130_fd_sc_hd__clkbuf_2 _22532_ (.A(\cpuregs_wrdata[8] ),
    .X(_19405_));
 sky130_fd_sc_hd__mux2_1 _22533_ (.A0(_19405_),
    .A1(\cpuregs[6][8] ),
    .S(_19400_),
    .X(_03704_));
 sky130_fd_sc_hd__clkbuf_2 _22534_ (.A(\cpuregs_wrdata[7] ),
    .X(_19406_));
 sky130_fd_sc_hd__buf_4 _22535_ (.A(_19377_),
    .X(_19407_));
 sky130_fd_sc_hd__mux2_1 _22536_ (.A0(_19406_),
    .A1(\cpuregs[6][7] ),
    .S(_19407_),
    .X(_03703_));
 sky130_fd_sc_hd__clkbuf_2 _22537_ (.A(\cpuregs_wrdata[6] ),
    .X(_19408_));
 sky130_fd_sc_hd__mux2_1 _22538_ (.A0(_19408_),
    .A1(\cpuregs[6][6] ),
    .S(_19407_),
    .X(_03702_));
 sky130_fd_sc_hd__clkbuf_2 _22539_ (.A(\cpuregs_wrdata[5] ),
    .X(_19409_));
 sky130_fd_sc_hd__mux2_1 _22540_ (.A0(_19409_),
    .A1(\cpuregs[6][5] ),
    .S(_19407_),
    .X(_03701_));
 sky130_fd_sc_hd__clkbuf_2 _22541_ (.A(\cpuregs_wrdata[4] ),
    .X(_19410_));
 sky130_fd_sc_hd__mux2_1 _22542_ (.A0(_19410_),
    .A1(\cpuregs[6][4] ),
    .S(_19407_),
    .X(_03700_));
 sky130_fd_sc_hd__clkbuf_2 _22543_ (.A(\cpuregs_wrdata[3] ),
    .X(_19411_));
 sky130_fd_sc_hd__mux2_1 _22544_ (.A0(_19411_),
    .A1(\cpuregs[6][3] ),
    .S(_19407_),
    .X(_03699_));
 sky130_fd_sc_hd__clkbuf_2 _22545_ (.A(\cpuregs_wrdata[2] ),
    .X(_19412_));
 sky130_fd_sc_hd__mux2_1 _22546_ (.A0(_19412_),
    .A1(\cpuregs[6][2] ),
    .S(_19407_),
    .X(_03698_));
 sky130_fd_sc_hd__clkbuf_2 _22547_ (.A(\cpuregs_wrdata[1] ),
    .X(_19413_));
 sky130_fd_sc_hd__mux2_1 _22548_ (.A0(_19413_),
    .A1(\cpuregs[6][1] ),
    .S(_19378_),
    .X(_03697_));
 sky130_fd_sc_hd__buf_1 _22549_ (.A(\cpuregs_wrdata[0] ),
    .X(_19414_));
 sky130_fd_sc_hd__mux2_1 _22550_ (.A0(_19414_),
    .A1(\cpuregs[6][0] ),
    .S(_19378_),
    .X(_03696_));
 sky130_fd_sc_hd__nor3_4 _22551_ (.A(_19365_),
    .B(\latched_rd[1] ),
    .C(_19372_),
    .Y(_19415_));
 sky130_fd_sc_hd__nand2_1 _22552_ (.A(_19367_),
    .B(\latched_rd[3] ),
    .Y(_19416_));
 sky130_vsdinv _22553_ (.A(_19416_),
    .Y(_19417_));
 sky130_fd_sc_hd__nand2_1 _22554_ (.A(_19415_),
    .B(_19417_),
    .Y(_19418_));
 sky130_fd_sc_hd__clkbuf_8 _22555_ (.A(_19418_),
    .X(_19419_));
 sky130_fd_sc_hd__buf_4 _22556_ (.A(_19419_),
    .X(_19420_));
 sky130_fd_sc_hd__mux2_1 _22557_ (.A0(_19363_),
    .A1(\cpuregs[9][31] ),
    .S(_19420_),
    .X(_03695_));
 sky130_fd_sc_hd__mux2_1 _22558_ (.A0(_19380_),
    .A1(\cpuregs[9][30] ),
    .S(_19420_),
    .X(_03694_));
 sky130_fd_sc_hd__mux2_1 _22559_ (.A0(_19381_),
    .A1(\cpuregs[9][29] ),
    .S(_19420_),
    .X(_03693_));
 sky130_fd_sc_hd__mux2_1 _22560_ (.A0(_19382_),
    .A1(\cpuregs[9][28] ),
    .S(_19420_),
    .X(_03692_));
 sky130_fd_sc_hd__mux2_1 _22561_ (.A0(_19383_),
    .A1(\cpuregs[9][27] ),
    .S(_19420_),
    .X(_03691_));
 sky130_fd_sc_hd__mux2_1 _22562_ (.A0(_19384_),
    .A1(\cpuregs[9][26] ),
    .S(_19420_),
    .X(_03690_));
 sky130_fd_sc_hd__buf_2 _22563_ (.A(_19419_),
    .X(_19421_));
 sky130_fd_sc_hd__mux2_1 _22564_ (.A0(_19385_),
    .A1(\cpuregs[9][25] ),
    .S(_19421_),
    .X(_03689_));
 sky130_fd_sc_hd__mux2_1 _22565_ (.A0(_19387_),
    .A1(\cpuregs[9][24] ),
    .S(_19421_),
    .X(_03688_));
 sky130_fd_sc_hd__mux2_1 _22566_ (.A0(_19388_),
    .A1(\cpuregs[9][23] ),
    .S(_19421_),
    .X(_03687_));
 sky130_fd_sc_hd__mux2_1 _22567_ (.A0(_19389_),
    .A1(\cpuregs[9][22] ),
    .S(_19421_),
    .X(_03686_));
 sky130_fd_sc_hd__mux2_1 _22568_ (.A0(_19390_),
    .A1(\cpuregs[9][21] ),
    .S(_19421_),
    .X(_03685_));
 sky130_fd_sc_hd__mux2_1 _22569_ (.A0(_19391_),
    .A1(\cpuregs[9][20] ),
    .S(_19421_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_4 _22570_ (.A(_19419_),
    .X(_19422_));
 sky130_fd_sc_hd__mux2_1 _22571_ (.A0(_19392_),
    .A1(\cpuregs[9][19] ),
    .S(_19422_),
    .X(_03683_));
 sky130_fd_sc_hd__mux2_1 _22572_ (.A0(_19394_),
    .A1(\cpuregs[9][18] ),
    .S(_19422_),
    .X(_03682_));
 sky130_fd_sc_hd__mux2_1 _22573_ (.A0(_19395_),
    .A1(\cpuregs[9][17] ),
    .S(_19422_),
    .X(_03681_));
 sky130_fd_sc_hd__mux2_1 _22574_ (.A0(_19396_),
    .A1(\cpuregs[9][16] ),
    .S(_19422_),
    .X(_03680_));
 sky130_fd_sc_hd__mux2_1 _22575_ (.A0(_19397_),
    .A1(\cpuregs[9][15] ),
    .S(_19422_),
    .X(_03679_));
 sky130_fd_sc_hd__mux2_1 _22576_ (.A0(_19398_),
    .A1(\cpuregs[9][14] ),
    .S(_19422_),
    .X(_03678_));
 sky130_fd_sc_hd__clkbuf_4 _22577_ (.A(_19419_),
    .X(_19423_));
 sky130_fd_sc_hd__mux2_1 _22578_ (.A0(_19399_),
    .A1(\cpuregs[9][13] ),
    .S(_19423_),
    .X(_03677_));
 sky130_fd_sc_hd__mux2_1 _22579_ (.A0(_19401_),
    .A1(\cpuregs[9][12] ),
    .S(_19423_),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_1 _22580_ (.A0(_19402_),
    .A1(\cpuregs[9][11] ),
    .S(_19423_),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_1 _22581_ (.A0(_19403_),
    .A1(\cpuregs[9][10] ),
    .S(_19423_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _22582_ (.A0(_19404_),
    .A1(\cpuregs[9][9] ),
    .S(_19423_),
    .X(_03673_));
 sky130_fd_sc_hd__mux2_1 _22583_ (.A0(_19405_),
    .A1(\cpuregs[9][8] ),
    .S(_19423_),
    .X(_03672_));
 sky130_fd_sc_hd__buf_4 _22584_ (.A(_19418_),
    .X(_19424_));
 sky130_fd_sc_hd__mux2_1 _22585_ (.A0(_19406_),
    .A1(\cpuregs[9][7] ),
    .S(_19424_),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _22586_ (.A0(_19408_),
    .A1(\cpuregs[9][6] ),
    .S(_19424_),
    .X(_03670_));
 sky130_fd_sc_hd__mux2_1 _22587_ (.A0(_19409_),
    .A1(\cpuregs[9][5] ),
    .S(_19424_),
    .X(_03669_));
 sky130_fd_sc_hd__mux2_1 _22588_ (.A0(_19410_),
    .A1(\cpuregs[9][4] ),
    .S(_19424_),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _22589_ (.A0(_19411_),
    .A1(\cpuregs[9][3] ),
    .S(_19424_),
    .X(_03667_));
 sky130_fd_sc_hd__mux2_1 _22590_ (.A0(_19412_),
    .A1(\cpuregs[9][2] ),
    .S(_19424_),
    .X(_03666_));
 sky130_fd_sc_hd__mux2_1 _22591_ (.A0(_19413_),
    .A1(\cpuregs[9][1] ),
    .S(_19419_),
    .X(_03665_));
 sky130_fd_sc_hd__mux2_1 _22592_ (.A0(_19414_),
    .A1(\cpuregs[9][0] ),
    .S(_19419_),
    .X(_03664_));
 sky130_fd_sc_hd__nor2_8 _22593_ (.A(_18310_),
    .B(_18498_),
    .Y(_19425_));
 sky130_fd_sc_hd__clkbuf_2 _22594_ (.A(_19425_),
    .X(_19426_));
 sky130_fd_sc_hd__clkbuf_4 _22595_ (.A(_19426_),
    .X(_19427_));
 sky130_fd_sc_hd__mux2_1 _22596_ (.A0(_18471_),
    .A1(_02467_),
    .S(_19427_),
    .X(_03663_));
 sky130_fd_sc_hd__buf_4 _22597_ (.A(net361),
    .X(_19428_));
 sky130_fd_sc_hd__mux2_1 _22598_ (.A0(_19428_),
    .A1(_02466_),
    .S(_19427_),
    .X(_03662_));
 sky130_fd_sc_hd__mux2_1 _22599_ (.A0(net359),
    .A1(_02464_),
    .S(_19427_),
    .X(_03661_));
 sky130_fd_sc_hd__mux2_1 _22600_ (.A0(net358),
    .A1(_02463_),
    .S(_19427_),
    .X(_03660_));
 sky130_fd_sc_hd__clkbuf_4 _22601_ (.A(net357),
    .X(_19429_));
 sky130_fd_sc_hd__mux2_1 _22602_ (.A0(_19429_),
    .A1(_02462_),
    .S(_19427_),
    .X(_03659_));
 sky130_fd_sc_hd__buf_2 _22603_ (.A(_19426_),
    .X(_19430_));
 sky130_fd_sc_hd__mux2_1 _22604_ (.A0(net356),
    .A1(_02461_),
    .S(_19430_),
    .X(_03658_));
 sky130_fd_sc_hd__mux2_1 _22605_ (.A0(net355),
    .A1(_02460_),
    .S(_19430_),
    .X(_03657_));
 sky130_fd_sc_hd__mux2_1 _22606_ (.A0(net354),
    .A1(_02459_),
    .S(_19430_),
    .X(_03656_));
 sky130_fd_sc_hd__clkbuf_4 _22607_ (.A(net353),
    .X(_19431_));
 sky130_fd_sc_hd__mux2_1 _22608_ (.A0(_19431_),
    .A1(_02458_),
    .S(_19430_),
    .X(_03655_));
 sky130_fd_sc_hd__buf_4 _22609_ (.A(net352),
    .X(_19432_));
 sky130_fd_sc_hd__mux2_1 _22610_ (.A0(_19432_),
    .A1(_02457_),
    .S(_19430_),
    .X(_03654_));
 sky130_fd_sc_hd__buf_4 _22611_ (.A(net351),
    .X(_19433_));
 sky130_fd_sc_hd__mux2_1 _22612_ (.A0(_19433_),
    .A1(_02456_),
    .S(_19430_),
    .X(_03653_));
 sky130_fd_sc_hd__clkbuf_4 _22613_ (.A(_19426_),
    .X(_19434_));
 sky130_fd_sc_hd__mux2_1 _22614_ (.A0(net350),
    .A1(_02455_),
    .S(_19434_),
    .X(_03652_));
 sky130_fd_sc_hd__mux2_1 _22615_ (.A0(net348),
    .A1(_02453_),
    .S(_19434_),
    .X(_03651_));
 sky130_fd_sc_hd__buf_4 _22616_ (.A(net347),
    .X(_19435_));
 sky130_fd_sc_hd__mux2_1 _22617_ (.A0(_19435_),
    .A1(_02452_),
    .S(_19434_),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_1 _22618_ (.A0(net346),
    .A1(_02451_),
    .S(_19434_),
    .X(_03649_));
 sky130_fd_sc_hd__buf_4 _22619_ (.A(net345),
    .X(_19436_));
 sky130_fd_sc_hd__mux2_1 _22620_ (.A0(_19436_),
    .A1(_02450_),
    .S(_19434_),
    .X(_03648_));
 sky130_fd_sc_hd__buf_4 _22621_ (.A(net344),
    .X(_19437_));
 sky130_fd_sc_hd__mux2_1 _22622_ (.A0(_19437_),
    .A1(_02449_),
    .S(_19434_),
    .X(_03647_));
 sky130_fd_sc_hd__buf_4 _22623_ (.A(net343),
    .X(_19438_));
 sky130_fd_sc_hd__buf_2 _22624_ (.A(_19425_),
    .X(_19439_));
 sky130_fd_sc_hd__mux2_1 _22625_ (.A0(_19438_),
    .A1(_02448_),
    .S(_19439_),
    .X(_03646_));
 sky130_fd_sc_hd__clkbuf_4 _22626_ (.A(net342),
    .X(_19440_));
 sky130_fd_sc_hd__mux2_1 _22627_ (.A0(_19440_),
    .A1(_02447_),
    .S(_19439_),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_4 _22628_ (.A(net341),
    .X(_19441_));
 sky130_fd_sc_hd__mux2_1 _22629_ (.A0(_19441_),
    .A1(_02446_),
    .S(_19439_),
    .X(_03644_));
 sky130_fd_sc_hd__clkbuf_4 _22630_ (.A(net340),
    .X(_19442_));
 sky130_fd_sc_hd__mux2_1 _22631_ (.A0(_19442_),
    .A1(_02445_),
    .S(_19439_),
    .X(_03643_));
 sky130_fd_sc_hd__buf_4 _22632_ (.A(net339),
    .X(_19443_));
 sky130_fd_sc_hd__mux2_1 _22633_ (.A0(_19443_),
    .A1(_02444_),
    .S(_19439_),
    .X(_03642_));
 sky130_fd_sc_hd__buf_4 _22634_ (.A(net369),
    .X(_19444_));
 sky130_fd_sc_hd__mux2_1 _22635_ (.A0(_19444_),
    .A1(_02474_),
    .S(_19439_),
    .X(_03641_));
 sky130_fd_sc_hd__buf_4 _22636_ (.A(net368),
    .X(_19445_));
 sky130_fd_sc_hd__buf_2 _22637_ (.A(_19425_),
    .X(_19446_));
 sky130_fd_sc_hd__mux2_1 _22638_ (.A0(_19445_),
    .A1(_02473_),
    .S(_19446_),
    .X(_03640_));
 sky130_fd_sc_hd__clkbuf_2 _22639_ (.A(net229),
    .X(_19447_));
 sky130_fd_sc_hd__mux2_1 _22640_ (.A0(net499),
    .A1(_02472_),
    .S(_19446_),
    .X(_03639_));
 sky130_fd_sc_hd__buf_6 _22641_ (.A(net228),
    .X(_19448_));
 sky130_fd_sc_hd__mux2_1 _22642_ (.A0(_19448_),
    .A1(_02471_),
    .S(_19446_),
    .X(_03638_));
 sky130_fd_sc_hd__buf_6 _22643_ (.A(net227),
    .X(_19449_));
 sky130_fd_sc_hd__mux2_1 _22644_ (.A0(_19449_),
    .A1(_02470_),
    .S(_19446_),
    .X(_03637_));
 sky130_fd_sc_hd__buf_6 _22645_ (.A(net226),
    .X(_19450_));
 sky130_fd_sc_hd__mux2_1 _22646_ (.A0(_19450_),
    .A1(_02469_),
    .S(_19446_),
    .X(_03636_));
 sky130_fd_sc_hd__buf_6 _22647_ (.A(net225),
    .X(_19451_));
 sky130_fd_sc_hd__mux2_1 _22648_ (.A0(_19451_),
    .A1(_02468_),
    .S(_19446_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_8 _22649_ (.A(net222),
    .X(_19452_));
 sky130_fd_sc_hd__mux2_1 _22650_ (.A0(_19452_),
    .A1(_02465_),
    .S(_19426_),
    .X(_03634_));
 sky130_fd_sc_hd__buf_4 _22651_ (.A(net211),
    .X(_19453_));
 sky130_fd_sc_hd__mux2_1 _22652_ (.A0(_19453_),
    .A1(_02454_),
    .S(_19426_),
    .X(_03633_));
 sky130_fd_sc_hd__buf_4 _22653_ (.A(net200),
    .X(_19454_));
 sky130_fd_sc_hd__mux2_1 _22654_ (.A0(_19454_),
    .A1(_02443_),
    .S(_19426_),
    .X(_03632_));
 sky130_fd_sc_hd__or3b_4 _22655_ (.A(_19366_),
    .B(_19372_),
    .C_N(_19376_),
    .X(_19455_));
 sky130_fd_sc_hd__clkbuf_8 _22656_ (.A(_19455_),
    .X(_19456_));
 sky130_fd_sc_hd__buf_4 _22657_ (.A(_19456_),
    .X(_19457_));
 sky130_fd_sc_hd__mux2_1 _22658_ (.A0(_19363_),
    .A1(\cpuregs[4][31] ),
    .S(_19457_),
    .X(_03631_));
 sky130_fd_sc_hd__mux2_1 _22659_ (.A0(_19380_),
    .A1(\cpuregs[4][30] ),
    .S(_19457_),
    .X(_03630_));
 sky130_fd_sc_hd__mux2_1 _22660_ (.A0(_19381_),
    .A1(\cpuregs[4][29] ),
    .S(_19457_),
    .X(_03629_));
 sky130_fd_sc_hd__mux2_1 _22661_ (.A0(_19382_),
    .A1(\cpuregs[4][28] ),
    .S(_19457_),
    .X(_03628_));
 sky130_fd_sc_hd__mux2_1 _22662_ (.A0(_19383_),
    .A1(\cpuregs[4][27] ),
    .S(_19457_),
    .X(_03627_));
 sky130_fd_sc_hd__mux2_1 _22663_ (.A0(_19384_),
    .A1(\cpuregs[4][26] ),
    .S(_19457_),
    .X(_03626_));
 sky130_fd_sc_hd__buf_2 _22664_ (.A(_19456_),
    .X(_19458_));
 sky130_fd_sc_hd__mux2_1 _22665_ (.A0(_19385_),
    .A1(\cpuregs[4][25] ),
    .S(_19458_),
    .X(_03625_));
 sky130_fd_sc_hd__mux2_1 _22666_ (.A0(_19387_),
    .A1(\cpuregs[4][24] ),
    .S(_19458_),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_1 _22667_ (.A0(_19388_),
    .A1(\cpuregs[4][23] ),
    .S(_19458_),
    .X(_03623_));
 sky130_fd_sc_hd__mux2_1 _22668_ (.A0(_19389_),
    .A1(\cpuregs[4][22] ),
    .S(_19458_),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_1 _22669_ (.A0(_19390_),
    .A1(\cpuregs[4][21] ),
    .S(_19458_),
    .X(_03621_));
 sky130_fd_sc_hd__mux2_1 _22670_ (.A0(_19391_),
    .A1(\cpuregs[4][20] ),
    .S(_19458_),
    .X(_03620_));
 sky130_fd_sc_hd__clkbuf_4 _22671_ (.A(_19456_),
    .X(_19459_));
 sky130_fd_sc_hd__mux2_1 _22672_ (.A0(_19392_),
    .A1(\cpuregs[4][19] ),
    .S(_19459_),
    .X(_03619_));
 sky130_fd_sc_hd__mux2_1 _22673_ (.A0(_19394_),
    .A1(\cpuregs[4][18] ),
    .S(_19459_),
    .X(_03618_));
 sky130_fd_sc_hd__mux2_1 _22674_ (.A0(_19395_),
    .A1(\cpuregs[4][17] ),
    .S(_19459_),
    .X(_03617_));
 sky130_fd_sc_hd__mux2_1 _22675_ (.A0(_19396_),
    .A1(\cpuregs[4][16] ),
    .S(_19459_),
    .X(_03616_));
 sky130_fd_sc_hd__mux2_1 _22676_ (.A0(_19397_),
    .A1(\cpuregs[4][15] ),
    .S(_19459_),
    .X(_03615_));
 sky130_fd_sc_hd__mux2_1 _22677_ (.A0(_19398_),
    .A1(\cpuregs[4][14] ),
    .S(_19459_),
    .X(_03614_));
 sky130_fd_sc_hd__clkbuf_4 _22678_ (.A(_19456_),
    .X(_19460_));
 sky130_fd_sc_hd__mux2_1 _22679_ (.A0(_19399_),
    .A1(\cpuregs[4][13] ),
    .S(_19460_),
    .X(_03613_));
 sky130_fd_sc_hd__mux2_1 _22680_ (.A0(_19401_),
    .A1(\cpuregs[4][12] ),
    .S(_19460_),
    .X(_03612_));
 sky130_fd_sc_hd__mux2_1 _22681_ (.A0(_19402_),
    .A1(\cpuregs[4][11] ),
    .S(_19460_),
    .X(_03611_));
 sky130_fd_sc_hd__mux2_1 _22682_ (.A0(_19403_),
    .A1(\cpuregs[4][10] ),
    .S(_19460_),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _22683_ (.A0(_19404_),
    .A1(\cpuregs[4][9] ),
    .S(_19460_),
    .X(_03609_));
 sky130_fd_sc_hd__mux2_1 _22684_ (.A0(_19405_),
    .A1(\cpuregs[4][8] ),
    .S(_19460_),
    .X(_03608_));
 sky130_fd_sc_hd__buf_4 _22685_ (.A(_19455_),
    .X(_19461_));
 sky130_fd_sc_hd__mux2_1 _22686_ (.A0(_19406_),
    .A1(\cpuregs[4][7] ),
    .S(_19461_),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _22687_ (.A0(_19408_),
    .A1(\cpuregs[4][6] ),
    .S(_19461_),
    .X(_03606_));
 sky130_fd_sc_hd__mux2_1 _22688_ (.A0(_19409_),
    .A1(\cpuregs[4][5] ),
    .S(_19461_),
    .X(_03605_));
 sky130_fd_sc_hd__mux2_1 _22689_ (.A0(_19410_),
    .A1(\cpuregs[4][4] ),
    .S(_19461_),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_1 _22690_ (.A0(_19411_),
    .A1(\cpuregs[4][3] ),
    .S(_19461_),
    .X(_03603_));
 sky130_fd_sc_hd__mux2_1 _22691_ (.A0(_19412_),
    .A1(\cpuregs[4][2] ),
    .S(_19461_),
    .X(_03602_));
 sky130_fd_sc_hd__mux2_1 _22692_ (.A0(_19413_),
    .A1(\cpuregs[4][1] ),
    .S(_19456_),
    .X(_03601_));
 sky130_fd_sc_hd__mux2_1 _22693_ (.A0(_19414_),
    .A1(\cpuregs[4][0] ),
    .S(_19456_),
    .X(_03600_));
 sky130_fd_sc_hd__nor2_4 _22694_ (.A(_19365_),
    .B(_19373_),
    .Y(_19462_));
 sky130_vsdinv _22695_ (.A(\latched_rd[2] ),
    .Y(_19463_));
 sky130_fd_sc_hd__and3_1 _22696_ (.A(_19463_),
    .B(_19368_),
    .C(\latched_rd[4] ),
    .X(_19464_));
 sky130_fd_sc_hd__nand2_1 _22697_ (.A(_19462_),
    .B(_19464_),
    .Y(_19465_));
 sky130_fd_sc_hd__buf_6 _22698_ (.A(_19465_),
    .X(_19466_));
 sky130_fd_sc_hd__clkbuf_4 _22699_ (.A(_19466_),
    .X(_19467_));
 sky130_fd_sc_hd__mux2_1 _22700_ (.A0(_19363_),
    .A1(\cpuregs[19][31] ),
    .S(_19467_),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_1 _22701_ (.A0(_19380_),
    .A1(\cpuregs[19][30] ),
    .S(_19467_),
    .X(_03598_));
 sky130_fd_sc_hd__mux2_1 _22702_ (.A0(_19381_),
    .A1(\cpuregs[19][29] ),
    .S(_19467_),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_1 _22703_ (.A0(_19382_),
    .A1(\cpuregs[19][28] ),
    .S(_19467_),
    .X(_03596_));
 sky130_fd_sc_hd__mux2_1 _22704_ (.A0(_19383_),
    .A1(\cpuregs[19][27] ),
    .S(_19467_),
    .X(_03595_));
 sky130_fd_sc_hd__mux2_1 _22705_ (.A0(_19384_),
    .A1(\cpuregs[19][26] ),
    .S(_19467_),
    .X(_03594_));
 sky130_fd_sc_hd__buf_2 _22706_ (.A(_19466_),
    .X(_19468_));
 sky130_fd_sc_hd__mux2_1 _22707_ (.A0(_19385_),
    .A1(\cpuregs[19][25] ),
    .S(_19468_),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_1 _22708_ (.A0(_19387_),
    .A1(\cpuregs[19][24] ),
    .S(_19468_),
    .X(_03592_));
 sky130_fd_sc_hd__mux2_1 _22709_ (.A0(_19388_),
    .A1(\cpuregs[19][23] ),
    .S(_19468_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_1 _22710_ (.A0(_19389_),
    .A1(\cpuregs[19][22] ),
    .S(_19468_),
    .X(_03590_));
 sky130_fd_sc_hd__mux2_1 _22711_ (.A0(_19390_),
    .A1(\cpuregs[19][21] ),
    .S(_19468_),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_1 _22712_ (.A0(_19391_),
    .A1(\cpuregs[19][20] ),
    .S(_19468_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_4 _22713_ (.A(_19466_),
    .X(_19469_));
 sky130_fd_sc_hd__mux2_1 _22714_ (.A0(_19392_),
    .A1(\cpuregs[19][19] ),
    .S(_19469_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _22715_ (.A0(_19394_),
    .A1(\cpuregs[19][18] ),
    .S(_19469_),
    .X(_03586_));
 sky130_fd_sc_hd__mux2_1 _22716_ (.A0(_19395_),
    .A1(\cpuregs[19][17] ),
    .S(_19469_),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_1 _22717_ (.A0(_19396_),
    .A1(\cpuregs[19][16] ),
    .S(_19469_),
    .X(_03584_));
 sky130_fd_sc_hd__mux2_1 _22718_ (.A0(_19397_),
    .A1(\cpuregs[19][15] ),
    .S(_19469_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _22719_ (.A0(_19398_),
    .A1(\cpuregs[19][14] ),
    .S(_19469_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_4 _22720_ (.A(_19466_),
    .X(_19470_));
 sky130_fd_sc_hd__mux2_1 _22721_ (.A0(_19399_),
    .A1(\cpuregs[19][13] ),
    .S(_19470_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_1 _22722_ (.A0(_19401_),
    .A1(\cpuregs[19][12] ),
    .S(_19470_),
    .X(_03580_));
 sky130_fd_sc_hd__mux2_1 _22723_ (.A0(_19402_),
    .A1(\cpuregs[19][11] ),
    .S(_19470_),
    .X(_03579_));
 sky130_fd_sc_hd__mux2_1 _22724_ (.A0(_19403_),
    .A1(\cpuregs[19][10] ),
    .S(_19470_),
    .X(_03578_));
 sky130_fd_sc_hd__mux2_1 _22725_ (.A0(_19404_),
    .A1(\cpuregs[19][9] ),
    .S(_19470_),
    .X(_03577_));
 sky130_fd_sc_hd__mux2_1 _22726_ (.A0(_19405_),
    .A1(\cpuregs[19][8] ),
    .S(_19470_),
    .X(_03576_));
 sky130_fd_sc_hd__clkbuf_4 _22727_ (.A(_19465_),
    .X(_19471_));
 sky130_fd_sc_hd__mux2_1 _22728_ (.A0(_19406_),
    .A1(\cpuregs[19][7] ),
    .S(_19471_),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_1 _22729_ (.A0(_19408_),
    .A1(\cpuregs[19][6] ),
    .S(_19471_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_1 _22730_ (.A0(_19409_),
    .A1(\cpuregs[19][5] ),
    .S(_19471_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _22731_ (.A0(_19410_),
    .A1(\cpuregs[19][4] ),
    .S(_19471_),
    .X(_03572_));
 sky130_fd_sc_hd__mux2_1 _22732_ (.A0(_19411_),
    .A1(\cpuregs[19][3] ),
    .S(_19471_),
    .X(_03571_));
 sky130_fd_sc_hd__mux2_1 _22733_ (.A0(_19412_),
    .A1(\cpuregs[19][2] ),
    .S(_19471_),
    .X(_03570_));
 sky130_fd_sc_hd__mux2_1 _22734_ (.A0(_19413_),
    .A1(\cpuregs[19][1] ),
    .S(_19466_),
    .X(_03569_));
 sky130_fd_sc_hd__mux2_1 _22735_ (.A0(_19414_),
    .A1(\cpuregs[19][0] ),
    .S(_19466_),
    .X(_03568_));
 sky130_fd_sc_hd__nor2_4 _22736_ (.A(_18309_),
    .B(_18317_),
    .Y(_19472_));
 sky130_fd_sc_hd__nand2_2 _22737_ (.A(_19472_),
    .B(_18630_),
    .Y(_19473_));
 sky130_fd_sc_hd__inv_4 _22738_ (.A(_19473_),
    .Y(net232));
 sky130_fd_sc_hd__nand2_2 _22739_ (.A(net232),
    .B(_18352_),
    .Y(_19474_));
 sky130_fd_sc_hd__buf_2 _22740_ (.A(_19474_),
    .X(_19475_));
 sky130_fd_sc_hd__buf_4 _22741_ (.A(_19475_),
    .X(_19476_));
 sky130_fd_sc_hd__mux2_1 _22742_ (.A0(net224),
    .A1(net262),
    .S(net421),
    .X(_03567_));
 sky130_fd_sc_hd__mux2_1 _22743_ (.A0(net223),
    .A1(net261),
    .S(net421),
    .X(_03566_));
 sky130_fd_sc_hd__mux2_1 _22744_ (.A0(net221),
    .A1(net259),
    .S(_19476_),
    .X(_03565_));
 sky130_fd_sc_hd__mux2_1 _22745_ (.A0(net220),
    .A1(net258),
    .S(net421),
    .X(_03564_));
 sky130_fd_sc_hd__mux2_1 _22746_ (.A0(net219),
    .A1(net257),
    .S(_19476_),
    .X(_03563_));
 sky130_fd_sc_hd__mux2_1 _22747_ (.A0(net218),
    .A1(net256),
    .S(net421),
    .X(_03562_));
 sky130_fd_sc_hd__buf_1 _22748_ (.A(_19475_),
    .X(_19477_));
 sky130_fd_sc_hd__mux2_1 _22749_ (.A0(net217),
    .A1(net255),
    .S(net420),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _22750_ (.A0(net216),
    .A1(net254),
    .S(net420),
    .X(_03560_));
 sky130_fd_sc_hd__mux2_1 _22751_ (.A0(net215),
    .A1(net253),
    .S(net420),
    .X(_03559_));
 sky130_fd_sc_hd__mux2_1 _22752_ (.A0(net214),
    .A1(net252),
    .S(net420),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_1 _22753_ (.A0(net213),
    .A1(net251),
    .S(net420),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_1 _22754_ (.A0(net212),
    .A1(net250),
    .S(net420),
    .X(_03556_));
 sky130_fd_sc_hd__buf_6 _22755_ (.A(_19475_),
    .X(_19478_));
 sky130_fd_sc_hd__mux2_1 _22756_ (.A0(net210),
    .A1(net248),
    .S(net419),
    .X(_03555_));
 sky130_fd_sc_hd__mux2_1 _22757_ (.A0(net209),
    .A1(net247),
    .S(_19478_),
    .X(_03554_));
 sky130_fd_sc_hd__mux2_1 _22758_ (.A0(net208),
    .A1(net246),
    .S(_19478_),
    .X(_03553_));
 sky130_fd_sc_hd__mux2_1 _22759_ (.A0(net207),
    .A1(net245),
    .S(_19478_),
    .X(_03552_));
 sky130_fd_sc_hd__mux2_1 _22760_ (.A0(net206),
    .A1(net244),
    .S(net419),
    .X(_03551_));
 sky130_fd_sc_hd__mux2_1 _22761_ (.A0(net205),
    .A1(net243),
    .S(net419),
    .X(_03550_));
 sky130_fd_sc_hd__buf_6 _22762_ (.A(_19475_),
    .X(_19479_));
 sky130_fd_sc_hd__mux2_1 _22763_ (.A0(net204),
    .A1(net242),
    .S(_19479_),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_1 _22764_ (.A0(net203),
    .A1(net241),
    .S(net418),
    .X(_03548_));
 sky130_fd_sc_hd__mux2_1 _22765_ (.A0(net202),
    .A1(net240),
    .S(net418),
    .X(_03547_));
 sky130_fd_sc_hd__mux2_1 _22766_ (.A0(net201),
    .A1(net239),
    .S(net418),
    .X(_03546_));
 sky130_fd_sc_hd__mux2_1 _22767_ (.A0(net231),
    .A1(net269),
    .S(_19479_),
    .X(_03545_));
 sky130_fd_sc_hd__mux2_1 _22768_ (.A0(net230),
    .A1(net268),
    .S(_19479_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_2 _22769_ (.A(_19474_),
    .X(_19480_));
 sky130_fd_sc_hd__mux2_1 _22770_ (.A0(net499),
    .A1(net267),
    .S(net423),
    .X(_03543_));
 sky130_fd_sc_hd__mux2_1 _22771_ (.A0(_19448_),
    .A1(net266),
    .S(net423),
    .X(_03542_));
 sky130_fd_sc_hd__mux2_1 _22772_ (.A0(_19449_),
    .A1(net265),
    .S(_19480_),
    .X(_03541_));
 sky130_fd_sc_hd__mux2_1 _22773_ (.A0(_19450_),
    .A1(net264),
    .S(net423),
    .X(_03540_));
 sky130_fd_sc_hd__mux2_1 _22774_ (.A0(_19451_),
    .A1(net263),
    .S(_19480_),
    .X(_03539_));
 sky130_fd_sc_hd__mux2_1 _22775_ (.A0(_19452_),
    .A1(net260),
    .S(net423),
    .X(_03538_));
 sky130_fd_sc_hd__mux2_1 _22776_ (.A0(_19453_),
    .A1(net249),
    .S(_19475_),
    .X(_03537_));
 sky130_fd_sc_hd__mux2_1 _22777_ (.A0(_19454_),
    .A1(net238),
    .S(_19475_),
    .X(_03536_));
 sky130_fd_sc_hd__nand2_1 _22778_ (.A(_19462_),
    .B(_19376_),
    .Y(_19481_));
 sky130_fd_sc_hd__clkbuf_8 _22779_ (.A(_19481_),
    .X(_19482_));
 sky130_fd_sc_hd__buf_4 _22780_ (.A(_19482_),
    .X(_19483_));
 sky130_fd_sc_hd__mux2_1 _22781_ (.A0(_19363_),
    .A1(\cpuregs[7][31] ),
    .S(_19483_),
    .X(_03535_));
 sky130_fd_sc_hd__mux2_1 _22782_ (.A0(_19380_),
    .A1(\cpuregs[7][30] ),
    .S(_19483_),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_1 _22783_ (.A0(_19381_),
    .A1(\cpuregs[7][29] ),
    .S(_19483_),
    .X(_03533_));
 sky130_fd_sc_hd__mux2_1 _22784_ (.A0(_19382_),
    .A1(\cpuregs[7][28] ),
    .S(_19483_),
    .X(_03532_));
 sky130_fd_sc_hd__mux2_1 _22785_ (.A0(_19383_),
    .A1(\cpuregs[7][27] ),
    .S(_19483_),
    .X(_03531_));
 sky130_fd_sc_hd__mux2_1 _22786_ (.A0(_19384_),
    .A1(\cpuregs[7][26] ),
    .S(_19483_),
    .X(_03530_));
 sky130_fd_sc_hd__buf_2 _22787_ (.A(_19482_),
    .X(_19484_));
 sky130_fd_sc_hd__mux2_1 _22788_ (.A0(_19385_),
    .A1(\cpuregs[7][25] ),
    .S(_19484_),
    .X(_03529_));
 sky130_fd_sc_hd__mux2_1 _22789_ (.A0(_19387_),
    .A1(\cpuregs[7][24] ),
    .S(_19484_),
    .X(_03528_));
 sky130_fd_sc_hd__mux2_1 _22790_ (.A0(_19388_),
    .A1(\cpuregs[7][23] ),
    .S(_19484_),
    .X(_03527_));
 sky130_fd_sc_hd__mux2_1 _22791_ (.A0(_19389_),
    .A1(\cpuregs[7][22] ),
    .S(_19484_),
    .X(_03526_));
 sky130_fd_sc_hd__mux2_1 _22792_ (.A0(_19390_),
    .A1(\cpuregs[7][21] ),
    .S(_19484_),
    .X(_03525_));
 sky130_fd_sc_hd__mux2_1 _22793_ (.A0(_19391_),
    .A1(\cpuregs[7][20] ),
    .S(_19484_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_4 _22794_ (.A(_19482_),
    .X(_19485_));
 sky130_fd_sc_hd__mux2_1 _22795_ (.A0(_19392_),
    .A1(\cpuregs[7][19] ),
    .S(_19485_),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_1 _22796_ (.A0(_19394_),
    .A1(\cpuregs[7][18] ),
    .S(_19485_),
    .X(_03522_));
 sky130_fd_sc_hd__mux2_1 _22797_ (.A0(_19395_),
    .A1(\cpuregs[7][17] ),
    .S(_19485_),
    .X(_03521_));
 sky130_fd_sc_hd__mux2_1 _22798_ (.A0(_19396_),
    .A1(\cpuregs[7][16] ),
    .S(_19485_),
    .X(_03520_));
 sky130_fd_sc_hd__mux2_1 _22799_ (.A0(_19397_),
    .A1(\cpuregs[7][15] ),
    .S(_19485_),
    .X(_03519_));
 sky130_fd_sc_hd__mux2_1 _22800_ (.A0(_19398_),
    .A1(\cpuregs[7][14] ),
    .S(_19485_),
    .X(_03518_));
 sky130_fd_sc_hd__buf_2 _22801_ (.A(_19482_),
    .X(_19486_));
 sky130_fd_sc_hd__mux2_1 _22802_ (.A0(_19399_),
    .A1(\cpuregs[7][13] ),
    .S(_19486_),
    .X(_03517_));
 sky130_fd_sc_hd__mux2_1 _22803_ (.A0(_19401_),
    .A1(\cpuregs[7][12] ),
    .S(_19486_),
    .X(_03516_));
 sky130_fd_sc_hd__mux2_1 _22804_ (.A0(_19402_),
    .A1(\cpuregs[7][11] ),
    .S(_19486_),
    .X(_03515_));
 sky130_fd_sc_hd__mux2_1 _22805_ (.A0(_19403_),
    .A1(\cpuregs[7][10] ),
    .S(_19486_),
    .X(_03514_));
 sky130_fd_sc_hd__mux2_1 _22806_ (.A0(_19404_),
    .A1(\cpuregs[7][9] ),
    .S(_19486_),
    .X(_03513_));
 sky130_fd_sc_hd__mux2_1 _22807_ (.A0(_19405_),
    .A1(\cpuregs[7][8] ),
    .S(_19486_),
    .X(_03512_));
 sky130_fd_sc_hd__buf_4 _22808_ (.A(_19481_),
    .X(_19487_));
 sky130_fd_sc_hd__mux2_1 _22809_ (.A0(_19406_),
    .A1(\cpuregs[7][7] ),
    .S(_19487_),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_1 _22810_ (.A0(_19408_),
    .A1(\cpuregs[7][6] ),
    .S(_19487_),
    .X(_03510_));
 sky130_fd_sc_hd__mux2_1 _22811_ (.A0(_19409_),
    .A1(\cpuregs[7][5] ),
    .S(_19487_),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_1 _22812_ (.A0(_19410_),
    .A1(\cpuregs[7][4] ),
    .S(_19487_),
    .X(_03508_));
 sky130_fd_sc_hd__mux2_1 _22813_ (.A0(_19411_),
    .A1(\cpuregs[7][3] ),
    .S(_19487_),
    .X(_03507_));
 sky130_fd_sc_hd__mux2_1 _22814_ (.A0(_19412_),
    .A1(\cpuregs[7][2] ),
    .S(_19487_),
    .X(_03506_));
 sky130_fd_sc_hd__mux2_1 _22815_ (.A0(_19413_),
    .A1(\cpuregs[7][1] ),
    .S(_19482_),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_1 _22816_ (.A0(_19414_),
    .A1(\cpuregs[7][0] ),
    .S(_19482_),
    .X(_03504_));
 sky130_fd_sc_hd__nor2_1 _22817_ (.A(_00331_),
    .B(_18310_),
    .Y(_19488_));
 sky130_fd_sc_hd__nand2_1 _22818_ (.A(_18540_),
    .B(_18481_),
    .Y(_19489_));
 sky130_fd_sc_hd__o211a_1 _22819_ (.A1(instr_setq),
    .A2(_19090_),
    .B1(_19488_),
    .C1(_19489_),
    .X(_19490_));
 sky130_fd_sc_hd__mux2_1 _22820_ (.A0(\latched_rd[4] ),
    .A1(_20891_),
    .S(_19490_),
    .X(_03503_));
 sky130_fd_sc_hd__and3_1 _22821_ (.A(_19375_),
    .B(\latched_rd[2] ),
    .C(\latched_rd[3] ),
    .X(_19491_));
 sky130_fd_sc_hd__nand2_1 _22822_ (.A(_19462_),
    .B(_19491_),
    .Y(_19492_));
 sky130_fd_sc_hd__clkbuf_8 _22823_ (.A(_19492_),
    .X(_19493_));
 sky130_fd_sc_hd__clkbuf_4 _22824_ (.A(_19493_),
    .X(_19494_));
 sky130_fd_sc_hd__mux2_1 _22825_ (.A0(_19363_),
    .A1(\cpuregs[15][31] ),
    .S(_19494_),
    .X(_03502_));
 sky130_fd_sc_hd__mux2_1 _22826_ (.A0(_19380_),
    .A1(\cpuregs[15][30] ),
    .S(_19494_),
    .X(_03501_));
 sky130_fd_sc_hd__mux2_1 _22827_ (.A0(_19381_),
    .A1(\cpuregs[15][29] ),
    .S(_19494_),
    .X(_03500_));
 sky130_fd_sc_hd__mux2_1 _22828_ (.A0(_19382_),
    .A1(\cpuregs[15][28] ),
    .S(_19494_),
    .X(_03499_));
 sky130_fd_sc_hd__mux2_1 _22829_ (.A0(_19383_),
    .A1(\cpuregs[15][27] ),
    .S(_19494_),
    .X(_03498_));
 sky130_fd_sc_hd__mux2_1 _22830_ (.A0(_19384_),
    .A1(\cpuregs[15][26] ),
    .S(_19494_),
    .X(_03497_));
 sky130_fd_sc_hd__buf_2 _22831_ (.A(_19493_),
    .X(_19495_));
 sky130_fd_sc_hd__mux2_1 _22832_ (.A0(_19385_),
    .A1(\cpuregs[15][25] ),
    .S(_19495_),
    .X(_03496_));
 sky130_fd_sc_hd__mux2_1 _22833_ (.A0(_19387_),
    .A1(\cpuregs[15][24] ),
    .S(_19495_),
    .X(_03495_));
 sky130_fd_sc_hd__mux2_1 _22834_ (.A0(_19388_),
    .A1(\cpuregs[15][23] ),
    .S(_19495_),
    .X(_03494_));
 sky130_fd_sc_hd__mux2_1 _22835_ (.A0(_19389_),
    .A1(\cpuregs[15][22] ),
    .S(_19495_),
    .X(_03493_));
 sky130_fd_sc_hd__mux2_1 _22836_ (.A0(_19390_),
    .A1(\cpuregs[15][21] ),
    .S(_19495_),
    .X(_03492_));
 sky130_fd_sc_hd__mux2_1 _22837_ (.A0(_19391_),
    .A1(\cpuregs[15][20] ),
    .S(_19495_),
    .X(_03491_));
 sky130_fd_sc_hd__buf_2 _22838_ (.A(_19493_),
    .X(_19496_));
 sky130_fd_sc_hd__mux2_1 _22839_ (.A0(_19392_),
    .A1(\cpuregs[15][19] ),
    .S(_19496_),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_1 _22840_ (.A0(_19394_),
    .A1(\cpuregs[15][18] ),
    .S(_19496_),
    .X(_03489_));
 sky130_fd_sc_hd__mux2_1 _22841_ (.A0(_19395_),
    .A1(\cpuregs[15][17] ),
    .S(_19496_),
    .X(_03488_));
 sky130_fd_sc_hd__mux2_1 _22842_ (.A0(_19396_),
    .A1(\cpuregs[15][16] ),
    .S(_19496_),
    .X(_03487_));
 sky130_fd_sc_hd__mux2_1 _22843_ (.A0(_19397_),
    .A1(\cpuregs[15][15] ),
    .S(_19496_),
    .X(_03486_));
 sky130_fd_sc_hd__mux2_1 _22844_ (.A0(_19398_),
    .A1(\cpuregs[15][14] ),
    .S(_19496_),
    .X(_03485_));
 sky130_fd_sc_hd__buf_2 _22845_ (.A(_19493_),
    .X(_19497_));
 sky130_fd_sc_hd__mux2_1 _22846_ (.A0(_19399_),
    .A1(\cpuregs[15][13] ),
    .S(_19497_),
    .X(_03484_));
 sky130_fd_sc_hd__mux2_1 _22847_ (.A0(_19401_),
    .A1(\cpuregs[15][12] ),
    .S(_19497_),
    .X(_03483_));
 sky130_fd_sc_hd__mux2_1 _22848_ (.A0(_19402_),
    .A1(\cpuregs[15][11] ),
    .S(_19497_),
    .X(_03482_));
 sky130_fd_sc_hd__mux2_1 _22849_ (.A0(_19403_),
    .A1(\cpuregs[15][10] ),
    .S(_19497_),
    .X(_03481_));
 sky130_fd_sc_hd__mux2_1 _22850_ (.A0(_19404_),
    .A1(\cpuregs[15][9] ),
    .S(_19497_),
    .X(_03480_));
 sky130_fd_sc_hd__mux2_1 _22851_ (.A0(_19405_),
    .A1(\cpuregs[15][8] ),
    .S(_19497_),
    .X(_03479_));
 sky130_fd_sc_hd__clkbuf_4 _22852_ (.A(_19492_),
    .X(_19498_));
 sky130_fd_sc_hd__mux2_1 _22853_ (.A0(_19406_),
    .A1(\cpuregs[15][7] ),
    .S(_19498_),
    .X(_03478_));
 sky130_fd_sc_hd__mux2_1 _22854_ (.A0(_19408_),
    .A1(\cpuregs[15][6] ),
    .S(_19498_),
    .X(_03477_));
 sky130_fd_sc_hd__mux2_1 _22855_ (.A0(_19409_),
    .A1(\cpuregs[15][5] ),
    .S(_19498_),
    .X(_03476_));
 sky130_fd_sc_hd__mux2_1 _22856_ (.A0(_19410_),
    .A1(\cpuregs[15][4] ),
    .S(_19498_),
    .X(_03475_));
 sky130_fd_sc_hd__mux2_1 _22857_ (.A0(_19411_),
    .A1(\cpuregs[15][3] ),
    .S(_19498_),
    .X(_03474_));
 sky130_fd_sc_hd__mux2_1 _22858_ (.A0(_19412_),
    .A1(\cpuregs[15][2] ),
    .S(_19498_),
    .X(_03473_));
 sky130_fd_sc_hd__mux2_1 _22859_ (.A0(_19413_),
    .A1(\cpuregs[15][1] ),
    .S(_19493_),
    .X(_03472_));
 sky130_fd_sc_hd__mux2_1 _22860_ (.A0(_19414_),
    .A1(\cpuregs[15][0] ),
    .S(_19493_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_2 _22861_ (.A(\cpuregs_wrdata[31] ),
    .X(_19499_));
 sky130_fd_sc_hd__nand2_1 _22862_ (.A(_19462_),
    .B(_19417_),
    .Y(_19500_));
 sky130_fd_sc_hd__buf_6 _22863_ (.A(_19500_),
    .X(_19501_));
 sky130_fd_sc_hd__clkbuf_4 _22864_ (.A(_19501_),
    .X(_19502_));
 sky130_fd_sc_hd__mux2_1 _22865_ (.A0(_19499_),
    .A1(\cpuregs[11][31] ),
    .S(_19502_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_2 _22866_ (.A(\cpuregs_wrdata[30] ),
    .X(_19503_));
 sky130_fd_sc_hd__mux2_1 _22867_ (.A0(_19503_),
    .A1(\cpuregs[11][30] ),
    .S(_19502_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_2 _22868_ (.A(\cpuregs_wrdata[29] ),
    .X(_19504_));
 sky130_fd_sc_hd__mux2_1 _22869_ (.A0(_19504_),
    .A1(\cpuregs[11][29] ),
    .S(_19502_),
    .X(_03468_));
 sky130_fd_sc_hd__clkbuf_2 _22870_ (.A(\cpuregs_wrdata[28] ),
    .X(_19505_));
 sky130_fd_sc_hd__mux2_1 _22871_ (.A0(_19505_),
    .A1(\cpuregs[11][28] ),
    .S(_19502_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_2 _22872_ (.A(\cpuregs_wrdata[27] ),
    .X(_19506_));
 sky130_fd_sc_hd__mux2_1 _22873_ (.A0(_19506_),
    .A1(\cpuregs[11][27] ),
    .S(_19502_),
    .X(_03466_));
 sky130_fd_sc_hd__clkbuf_2 _22874_ (.A(\cpuregs_wrdata[26] ),
    .X(_19507_));
 sky130_fd_sc_hd__mux2_1 _22875_ (.A0(_19507_),
    .A1(\cpuregs[11][26] ),
    .S(_19502_),
    .X(_03465_));
 sky130_fd_sc_hd__clkbuf_2 _22876_ (.A(\cpuregs_wrdata[25] ),
    .X(_19508_));
 sky130_fd_sc_hd__buf_2 _22877_ (.A(_19501_),
    .X(_19509_));
 sky130_fd_sc_hd__mux2_1 _22878_ (.A0(_19508_),
    .A1(\cpuregs[11][25] ),
    .S(_19509_),
    .X(_03464_));
 sky130_fd_sc_hd__clkbuf_2 _22879_ (.A(\cpuregs_wrdata[24] ),
    .X(_19510_));
 sky130_fd_sc_hd__mux2_1 _22880_ (.A0(_19510_),
    .A1(\cpuregs[11][24] ),
    .S(_19509_),
    .X(_03463_));
 sky130_fd_sc_hd__clkbuf_2 _22881_ (.A(\cpuregs_wrdata[23] ),
    .X(_19511_));
 sky130_fd_sc_hd__mux2_1 _22882_ (.A0(_19511_),
    .A1(\cpuregs[11][23] ),
    .S(_19509_),
    .X(_03462_));
 sky130_fd_sc_hd__clkbuf_2 _22883_ (.A(\cpuregs_wrdata[22] ),
    .X(_19512_));
 sky130_fd_sc_hd__mux2_1 _22884_ (.A0(_19512_),
    .A1(\cpuregs[11][22] ),
    .S(_19509_),
    .X(_03461_));
 sky130_fd_sc_hd__clkbuf_2 _22885_ (.A(\cpuregs_wrdata[21] ),
    .X(_19513_));
 sky130_fd_sc_hd__mux2_1 _22886_ (.A0(_19513_),
    .A1(\cpuregs[11][21] ),
    .S(_19509_),
    .X(_03460_));
 sky130_fd_sc_hd__clkbuf_2 _22887_ (.A(\cpuregs_wrdata[20] ),
    .X(_19514_));
 sky130_fd_sc_hd__mux2_1 _22888_ (.A0(_19514_),
    .A1(\cpuregs[11][20] ),
    .S(_19509_),
    .X(_03459_));
 sky130_fd_sc_hd__clkbuf_2 _22889_ (.A(\cpuregs_wrdata[19] ),
    .X(_19515_));
 sky130_fd_sc_hd__clkbuf_4 _22890_ (.A(_19501_),
    .X(_19516_));
 sky130_fd_sc_hd__mux2_1 _22891_ (.A0(_19515_),
    .A1(\cpuregs[11][19] ),
    .S(_19516_),
    .X(_03458_));
 sky130_fd_sc_hd__clkbuf_2 _22892_ (.A(\cpuregs_wrdata[18] ),
    .X(_19517_));
 sky130_fd_sc_hd__mux2_1 _22893_ (.A0(_19517_),
    .A1(\cpuregs[11][18] ),
    .S(_19516_),
    .X(_03457_));
 sky130_fd_sc_hd__clkbuf_2 _22894_ (.A(\cpuregs_wrdata[17] ),
    .X(_19518_));
 sky130_fd_sc_hd__mux2_1 _22895_ (.A0(_19518_),
    .A1(\cpuregs[11][17] ),
    .S(_19516_),
    .X(_03456_));
 sky130_fd_sc_hd__clkbuf_2 _22896_ (.A(\cpuregs_wrdata[16] ),
    .X(_19519_));
 sky130_fd_sc_hd__mux2_1 _22897_ (.A0(_19519_),
    .A1(\cpuregs[11][16] ),
    .S(_19516_),
    .X(_03455_));
 sky130_fd_sc_hd__clkbuf_2 _22898_ (.A(\cpuregs_wrdata[15] ),
    .X(_19520_));
 sky130_fd_sc_hd__mux2_1 _22899_ (.A0(_19520_),
    .A1(\cpuregs[11][15] ),
    .S(_19516_),
    .X(_03454_));
 sky130_fd_sc_hd__clkbuf_2 _22900_ (.A(\cpuregs_wrdata[14] ),
    .X(_19521_));
 sky130_fd_sc_hd__mux2_1 _22901_ (.A0(_19521_),
    .A1(\cpuregs[11][14] ),
    .S(_19516_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_2 _22902_ (.A(\cpuregs_wrdata[13] ),
    .X(_19522_));
 sky130_fd_sc_hd__buf_2 _22903_ (.A(_19501_),
    .X(_19523_));
 sky130_fd_sc_hd__mux2_1 _22904_ (.A0(_19522_),
    .A1(\cpuregs[11][13] ),
    .S(_19523_),
    .X(_03452_));
 sky130_fd_sc_hd__clkbuf_2 _22905_ (.A(\cpuregs_wrdata[12] ),
    .X(_19524_));
 sky130_fd_sc_hd__mux2_1 _22906_ (.A0(_19524_),
    .A1(\cpuregs[11][12] ),
    .S(_19523_),
    .X(_03451_));
 sky130_fd_sc_hd__clkbuf_2 _22907_ (.A(\cpuregs_wrdata[11] ),
    .X(_19525_));
 sky130_fd_sc_hd__mux2_1 _22908_ (.A0(_19525_),
    .A1(\cpuregs[11][11] ),
    .S(_19523_),
    .X(_03450_));
 sky130_fd_sc_hd__clkbuf_2 _22909_ (.A(\cpuregs_wrdata[10] ),
    .X(_19526_));
 sky130_fd_sc_hd__mux2_1 _22910_ (.A0(_19526_),
    .A1(\cpuregs[11][10] ),
    .S(_19523_),
    .X(_03449_));
 sky130_fd_sc_hd__clkbuf_2 _22911_ (.A(\cpuregs_wrdata[9] ),
    .X(_19527_));
 sky130_fd_sc_hd__mux2_1 _22912_ (.A0(_19527_),
    .A1(\cpuregs[11][9] ),
    .S(_19523_),
    .X(_03448_));
 sky130_fd_sc_hd__clkbuf_2 _22913_ (.A(\cpuregs_wrdata[8] ),
    .X(_19528_));
 sky130_fd_sc_hd__mux2_1 _22914_ (.A0(_19528_),
    .A1(\cpuregs[11][8] ),
    .S(_19523_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_2 _22915_ (.A(\cpuregs_wrdata[7] ),
    .X(_19529_));
 sky130_fd_sc_hd__clkbuf_4 _22916_ (.A(_19500_),
    .X(_19530_));
 sky130_fd_sc_hd__mux2_1 _22917_ (.A0(_19529_),
    .A1(\cpuregs[11][7] ),
    .S(_19530_),
    .X(_03446_));
 sky130_fd_sc_hd__clkbuf_2 _22918_ (.A(\cpuregs_wrdata[6] ),
    .X(_19531_));
 sky130_fd_sc_hd__mux2_1 _22919_ (.A0(_19531_),
    .A1(\cpuregs[11][6] ),
    .S(_19530_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_2 _22920_ (.A(\cpuregs_wrdata[5] ),
    .X(_19532_));
 sky130_fd_sc_hd__mux2_1 _22921_ (.A0(_19532_),
    .A1(\cpuregs[11][5] ),
    .S(_19530_),
    .X(_03444_));
 sky130_fd_sc_hd__clkbuf_2 _22922_ (.A(\cpuregs_wrdata[4] ),
    .X(_19533_));
 sky130_fd_sc_hd__mux2_1 _22923_ (.A0(_19533_),
    .A1(\cpuregs[11][4] ),
    .S(_19530_),
    .X(_03443_));
 sky130_fd_sc_hd__buf_1 _22924_ (.A(\cpuregs_wrdata[3] ),
    .X(_19534_));
 sky130_fd_sc_hd__mux2_1 _22925_ (.A0(_19534_),
    .A1(\cpuregs[11][3] ),
    .S(_19530_),
    .X(_03442_));
 sky130_fd_sc_hd__clkbuf_2 _22926_ (.A(\cpuregs_wrdata[2] ),
    .X(_19535_));
 sky130_fd_sc_hd__mux2_1 _22927_ (.A0(_19535_),
    .A1(\cpuregs[11][2] ),
    .S(_19530_),
    .X(_03441_));
 sky130_fd_sc_hd__clkbuf_2 _22928_ (.A(\cpuregs_wrdata[1] ),
    .X(_19536_));
 sky130_fd_sc_hd__mux2_1 _22929_ (.A0(_19536_),
    .A1(\cpuregs[11][1] ),
    .S(_19501_),
    .X(_03440_));
 sky130_fd_sc_hd__clkbuf_2 _22930_ (.A(\cpuregs_wrdata[0] ),
    .X(_19537_));
 sky130_fd_sc_hd__mux2_1 _22931_ (.A0(_19537_),
    .A1(\cpuregs[11][0] ),
    .S(_19501_),
    .X(_03439_));
 sky130_vsdinv _22932_ (.A(_19369_),
    .Y(_19538_));
 sky130_fd_sc_hd__nand2_2 _22933_ (.A(_19462_),
    .B(_19538_),
    .Y(_19539_));
 sky130_fd_sc_hd__buf_8 _22934_ (.A(_19539_),
    .X(_19540_));
 sky130_fd_sc_hd__clkbuf_4 _22935_ (.A(_19540_),
    .X(_19541_));
 sky130_fd_sc_hd__mux2_1 _22936_ (.A0(_19499_),
    .A1(\cpuregs[3][31] ),
    .S(_19541_),
    .X(_03438_));
 sky130_fd_sc_hd__mux2_1 _22937_ (.A0(_19503_),
    .A1(\cpuregs[3][30] ),
    .S(_19541_),
    .X(_03437_));
 sky130_fd_sc_hd__mux2_1 _22938_ (.A0(_19504_),
    .A1(\cpuregs[3][29] ),
    .S(_19541_),
    .X(_03436_));
 sky130_fd_sc_hd__mux2_1 _22939_ (.A0(_19505_),
    .A1(\cpuregs[3][28] ),
    .S(_19541_),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _22940_ (.A0(_19506_),
    .A1(\cpuregs[3][27] ),
    .S(_19541_),
    .X(_03434_));
 sky130_fd_sc_hd__mux2_1 _22941_ (.A0(_19507_),
    .A1(\cpuregs[3][26] ),
    .S(_19541_),
    .X(_03433_));
 sky130_fd_sc_hd__buf_2 _22942_ (.A(_19540_),
    .X(_19542_));
 sky130_fd_sc_hd__mux2_1 _22943_ (.A0(_19508_),
    .A1(\cpuregs[3][25] ),
    .S(_19542_),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_1 _22944_ (.A0(_19510_),
    .A1(\cpuregs[3][24] ),
    .S(_19542_),
    .X(_03431_));
 sky130_fd_sc_hd__mux2_1 _22945_ (.A0(_19511_),
    .A1(\cpuregs[3][23] ),
    .S(_19542_),
    .X(_03430_));
 sky130_fd_sc_hd__mux2_1 _22946_ (.A0(_19512_),
    .A1(\cpuregs[3][22] ),
    .S(_19542_),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_1 _22947_ (.A0(_19513_),
    .A1(\cpuregs[3][21] ),
    .S(_19542_),
    .X(_03428_));
 sky130_fd_sc_hd__mux2_1 _22948_ (.A0(_19514_),
    .A1(\cpuregs[3][20] ),
    .S(_19542_),
    .X(_03427_));
 sky130_fd_sc_hd__clkbuf_4 _22949_ (.A(_19540_),
    .X(_19543_));
 sky130_fd_sc_hd__mux2_1 _22950_ (.A0(_19515_),
    .A1(\cpuregs[3][19] ),
    .S(_19543_),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _22951_ (.A0(_19517_),
    .A1(\cpuregs[3][18] ),
    .S(_19543_),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_1 _22952_ (.A0(_19518_),
    .A1(\cpuregs[3][17] ),
    .S(_19543_),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_1 _22953_ (.A0(_19519_),
    .A1(\cpuregs[3][16] ),
    .S(_19543_),
    .X(_03423_));
 sky130_fd_sc_hd__mux2_1 _22954_ (.A0(_19520_),
    .A1(\cpuregs[3][15] ),
    .S(_19543_),
    .X(_03422_));
 sky130_fd_sc_hd__mux2_1 _22955_ (.A0(_19521_),
    .A1(\cpuregs[3][14] ),
    .S(_19543_),
    .X(_03421_));
 sky130_fd_sc_hd__buf_2 _22956_ (.A(_19540_),
    .X(_19544_));
 sky130_fd_sc_hd__mux2_1 _22957_ (.A0(_19522_),
    .A1(\cpuregs[3][13] ),
    .S(_19544_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _22958_ (.A0(_19524_),
    .A1(\cpuregs[3][12] ),
    .S(_19544_),
    .X(_03419_));
 sky130_fd_sc_hd__mux2_1 _22959_ (.A0(_19525_),
    .A1(\cpuregs[3][11] ),
    .S(_19544_),
    .X(_03418_));
 sky130_fd_sc_hd__mux2_1 _22960_ (.A0(_19526_),
    .A1(\cpuregs[3][10] ),
    .S(_19544_),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_1 _22961_ (.A0(_19527_),
    .A1(\cpuregs[3][9] ),
    .S(_19544_),
    .X(_03416_));
 sky130_fd_sc_hd__mux2_1 _22962_ (.A0(_19528_),
    .A1(\cpuregs[3][8] ),
    .S(_19544_),
    .X(_03415_));
 sky130_fd_sc_hd__buf_4 _22963_ (.A(_19539_),
    .X(_19545_));
 sky130_fd_sc_hd__mux2_1 _22964_ (.A0(_19529_),
    .A1(\cpuregs[3][7] ),
    .S(_19545_),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _22965_ (.A0(_19531_),
    .A1(\cpuregs[3][6] ),
    .S(_19545_),
    .X(_03413_));
 sky130_fd_sc_hd__mux2_1 _22966_ (.A0(_19532_),
    .A1(\cpuregs[3][5] ),
    .S(_19545_),
    .X(_03412_));
 sky130_fd_sc_hd__mux2_1 _22967_ (.A0(_19533_),
    .A1(\cpuregs[3][4] ),
    .S(_19545_),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_1 _22968_ (.A0(_19534_),
    .A1(\cpuregs[3][3] ),
    .S(_19545_),
    .X(_03410_));
 sky130_fd_sc_hd__mux2_1 _22969_ (.A0(_19535_),
    .A1(\cpuregs[3][2] ),
    .S(_19545_),
    .X(_03409_));
 sky130_fd_sc_hd__mux2_1 _22970_ (.A0(_19536_),
    .A1(\cpuregs[3][1] ),
    .S(_19540_),
    .X(_03408_));
 sky130_fd_sc_hd__mux2_1 _22971_ (.A0(_19537_),
    .A1(\cpuregs[3][0] ),
    .S(_19540_),
    .X(_03407_));
 sky130_fd_sc_hd__nand2_1 _22972_ (.A(_19415_),
    .B(_19538_),
    .Y(_19546_));
 sky130_fd_sc_hd__buf_8 _22973_ (.A(_19546_),
    .X(_19547_));
 sky130_fd_sc_hd__clkbuf_4 _22974_ (.A(_19547_),
    .X(_19548_));
 sky130_fd_sc_hd__mux2_1 _22975_ (.A0(_19499_),
    .A1(\cpuregs[1][31] ),
    .S(_19548_),
    .X(_03406_));
 sky130_fd_sc_hd__mux2_1 _22976_ (.A0(_19503_),
    .A1(\cpuregs[1][30] ),
    .S(_19548_),
    .X(_03405_));
 sky130_fd_sc_hd__mux2_1 _22977_ (.A0(_19504_),
    .A1(\cpuregs[1][29] ),
    .S(_19548_),
    .X(_03404_));
 sky130_fd_sc_hd__mux2_1 _22978_ (.A0(_19505_),
    .A1(\cpuregs[1][28] ),
    .S(_19548_),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_1 _22979_ (.A0(_19506_),
    .A1(\cpuregs[1][27] ),
    .S(_19548_),
    .X(_03402_));
 sky130_fd_sc_hd__mux2_1 _22980_ (.A0(_19507_),
    .A1(\cpuregs[1][26] ),
    .S(_19548_),
    .X(_03401_));
 sky130_fd_sc_hd__buf_2 _22981_ (.A(_19547_),
    .X(_19549_));
 sky130_fd_sc_hd__mux2_1 _22982_ (.A0(_19508_),
    .A1(\cpuregs[1][25] ),
    .S(_19549_),
    .X(_03400_));
 sky130_fd_sc_hd__mux2_1 _22983_ (.A0(_19510_),
    .A1(\cpuregs[1][24] ),
    .S(_19549_),
    .X(_03399_));
 sky130_fd_sc_hd__mux2_1 _22984_ (.A0(_19511_),
    .A1(\cpuregs[1][23] ),
    .S(_19549_),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_1 _22985_ (.A0(_19512_),
    .A1(\cpuregs[1][22] ),
    .S(_19549_),
    .X(_03397_));
 sky130_fd_sc_hd__mux2_1 _22986_ (.A0(_19513_),
    .A1(\cpuregs[1][21] ),
    .S(_19549_),
    .X(_03396_));
 sky130_fd_sc_hd__mux2_1 _22987_ (.A0(_19514_),
    .A1(\cpuregs[1][20] ),
    .S(_19549_),
    .X(_03395_));
 sky130_fd_sc_hd__clkbuf_4 _22988_ (.A(_19547_),
    .X(_19550_));
 sky130_fd_sc_hd__mux2_1 _22989_ (.A0(_19515_),
    .A1(\cpuregs[1][19] ),
    .S(_19550_),
    .X(_03394_));
 sky130_fd_sc_hd__mux2_1 _22990_ (.A0(_19517_),
    .A1(\cpuregs[1][18] ),
    .S(_19550_),
    .X(_03393_));
 sky130_fd_sc_hd__mux2_1 _22991_ (.A0(_19518_),
    .A1(\cpuregs[1][17] ),
    .S(_19550_),
    .X(_03392_));
 sky130_fd_sc_hd__mux2_1 _22992_ (.A0(_19519_),
    .A1(\cpuregs[1][16] ),
    .S(_19550_),
    .X(_03391_));
 sky130_fd_sc_hd__mux2_1 _22993_ (.A0(_19520_),
    .A1(\cpuregs[1][15] ),
    .S(_19550_),
    .X(_03390_));
 sky130_fd_sc_hd__mux2_1 _22994_ (.A0(_19521_),
    .A1(\cpuregs[1][14] ),
    .S(_19550_),
    .X(_03389_));
 sky130_fd_sc_hd__buf_2 _22995_ (.A(_19547_),
    .X(_19551_));
 sky130_fd_sc_hd__mux2_1 _22996_ (.A0(_19522_),
    .A1(\cpuregs[1][13] ),
    .S(_19551_),
    .X(_03388_));
 sky130_fd_sc_hd__mux2_1 _22997_ (.A0(_19524_),
    .A1(\cpuregs[1][12] ),
    .S(_19551_),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _22998_ (.A0(_19525_),
    .A1(\cpuregs[1][11] ),
    .S(_19551_),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_1 _22999_ (.A0(_19526_),
    .A1(\cpuregs[1][10] ),
    .S(_19551_),
    .X(_03385_));
 sky130_fd_sc_hd__mux2_1 _23000_ (.A0(_19527_),
    .A1(\cpuregs[1][9] ),
    .S(_19551_),
    .X(_03384_));
 sky130_fd_sc_hd__mux2_1 _23001_ (.A0(_19528_),
    .A1(\cpuregs[1][8] ),
    .S(_19551_),
    .X(_03383_));
 sky130_fd_sc_hd__buf_4 _23002_ (.A(_19546_),
    .X(_19552_));
 sky130_fd_sc_hd__mux2_1 _23003_ (.A0(_19529_),
    .A1(\cpuregs[1][7] ),
    .S(_19552_),
    .X(_03382_));
 sky130_fd_sc_hd__mux2_1 _23004_ (.A0(_19531_),
    .A1(\cpuregs[1][6] ),
    .S(_19552_),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_1 _23005_ (.A0(_19532_),
    .A1(\cpuregs[1][5] ),
    .S(_19552_),
    .X(_03380_));
 sky130_fd_sc_hd__mux2_1 _23006_ (.A0(_19533_),
    .A1(\cpuregs[1][4] ),
    .S(_19552_),
    .X(_03379_));
 sky130_fd_sc_hd__mux2_1 _23007_ (.A0(_19534_),
    .A1(\cpuregs[1][3] ),
    .S(_19552_),
    .X(_03378_));
 sky130_fd_sc_hd__mux2_1 _23008_ (.A0(_19535_),
    .A1(\cpuregs[1][2] ),
    .S(_19552_),
    .X(_03377_));
 sky130_fd_sc_hd__mux2_1 _23009_ (.A0(_19536_),
    .A1(\cpuregs[1][1] ),
    .S(_19547_),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_1 _23010_ (.A0(_19537_),
    .A1(\cpuregs[1][0] ),
    .S(_19547_),
    .X(_03375_));
 sky130_fd_sc_hd__or3b_4 _23011_ (.A(_19366_),
    .B(_19372_),
    .C_N(_19491_),
    .X(_19553_));
 sky130_fd_sc_hd__buf_8 _23012_ (.A(_19553_),
    .X(_19554_));
 sky130_fd_sc_hd__clkbuf_4 _23013_ (.A(_19554_),
    .X(_19555_));
 sky130_fd_sc_hd__mux2_1 _23014_ (.A0(_19499_),
    .A1(\cpuregs[12][31] ),
    .S(_19555_),
    .X(_03374_));
 sky130_fd_sc_hd__mux2_1 _23015_ (.A0(_19503_),
    .A1(\cpuregs[12][30] ),
    .S(_19555_),
    .X(_03373_));
 sky130_fd_sc_hd__mux2_1 _23016_ (.A0(_19504_),
    .A1(\cpuregs[12][29] ),
    .S(_19555_),
    .X(_03372_));
 sky130_fd_sc_hd__mux2_1 _23017_ (.A0(_19505_),
    .A1(\cpuregs[12][28] ),
    .S(_19555_),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_1 _23018_ (.A0(_19506_),
    .A1(\cpuregs[12][27] ),
    .S(_19555_),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_1 _23019_ (.A0(_19507_),
    .A1(\cpuregs[12][26] ),
    .S(_19555_),
    .X(_03369_));
 sky130_fd_sc_hd__buf_2 _23020_ (.A(_19554_),
    .X(_19556_));
 sky130_fd_sc_hd__mux2_1 _23021_ (.A0(_19508_),
    .A1(\cpuregs[12][25] ),
    .S(_19556_),
    .X(_03368_));
 sky130_fd_sc_hd__mux2_1 _23022_ (.A0(_19510_),
    .A1(\cpuregs[12][24] ),
    .S(_19556_),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_1 _23023_ (.A0(_19511_),
    .A1(\cpuregs[12][23] ),
    .S(_19556_),
    .X(_03366_));
 sky130_fd_sc_hd__mux2_1 _23024_ (.A0(_19512_),
    .A1(\cpuregs[12][22] ),
    .S(_19556_),
    .X(_03365_));
 sky130_fd_sc_hd__mux2_1 _23025_ (.A0(_19513_),
    .A1(\cpuregs[12][21] ),
    .S(_19556_),
    .X(_03364_));
 sky130_fd_sc_hd__mux2_1 _23026_ (.A0(_19514_),
    .A1(\cpuregs[12][20] ),
    .S(_19556_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_4 _23027_ (.A(_19554_),
    .X(_19557_));
 sky130_fd_sc_hd__mux2_1 _23028_ (.A0(_19515_),
    .A1(\cpuregs[12][19] ),
    .S(_19557_),
    .X(_03362_));
 sky130_fd_sc_hd__mux2_1 _23029_ (.A0(_19517_),
    .A1(\cpuregs[12][18] ),
    .S(_19557_),
    .X(_03361_));
 sky130_fd_sc_hd__mux2_1 _23030_ (.A0(_19518_),
    .A1(\cpuregs[12][17] ),
    .S(_19557_),
    .X(_03360_));
 sky130_fd_sc_hd__mux2_1 _23031_ (.A0(_19519_),
    .A1(\cpuregs[12][16] ),
    .S(_19557_),
    .X(_03359_));
 sky130_fd_sc_hd__mux2_1 _23032_ (.A0(_19520_),
    .A1(\cpuregs[12][15] ),
    .S(_19557_),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_1 _23033_ (.A0(_19521_),
    .A1(\cpuregs[12][14] ),
    .S(_19557_),
    .X(_03357_));
 sky130_fd_sc_hd__buf_2 _23034_ (.A(_19554_),
    .X(_19558_));
 sky130_fd_sc_hd__mux2_1 _23035_ (.A0(_19522_),
    .A1(\cpuregs[12][13] ),
    .S(_19558_),
    .X(_03356_));
 sky130_fd_sc_hd__mux2_1 _23036_ (.A0(_19524_),
    .A1(\cpuregs[12][12] ),
    .S(_19558_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _23037_ (.A0(_19525_),
    .A1(\cpuregs[12][11] ),
    .S(_19558_),
    .X(_03354_));
 sky130_fd_sc_hd__mux2_1 _23038_ (.A0(_19526_),
    .A1(\cpuregs[12][10] ),
    .S(_19558_),
    .X(_03353_));
 sky130_fd_sc_hd__mux2_1 _23039_ (.A0(_19527_),
    .A1(\cpuregs[12][9] ),
    .S(_19558_),
    .X(_03352_));
 sky130_fd_sc_hd__mux2_1 _23040_ (.A0(_19528_),
    .A1(\cpuregs[12][8] ),
    .S(_19558_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_4 _23041_ (.A(_19553_),
    .X(_19559_));
 sky130_fd_sc_hd__mux2_1 _23042_ (.A0(_19529_),
    .A1(\cpuregs[12][7] ),
    .S(_19559_),
    .X(_03350_));
 sky130_fd_sc_hd__mux2_1 _23043_ (.A0(_19531_),
    .A1(\cpuregs[12][6] ),
    .S(_19559_),
    .X(_03349_));
 sky130_fd_sc_hd__mux2_1 _23044_ (.A0(_19532_),
    .A1(\cpuregs[12][5] ),
    .S(_19559_),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _23045_ (.A0(_19533_),
    .A1(\cpuregs[12][4] ),
    .S(_19559_),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_1 _23046_ (.A0(_19534_),
    .A1(\cpuregs[12][3] ),
    .S(_19559_),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_1 _23047_ (.A0(_19535_),
    .A1(\cpuregs[12][2] ),
    .S(_19559_),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _23048_ (.A0(_19536_),
    .A1(\cpuregs[12][1] ),
    .S(_19554_),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_1 _23049_ (.A0(_19537_),
    .A1(\cpuregs[12][0] ),
    .S(_19554_),
    .X(_03343_));
 sky130_fd_sc_hd__or3_2 _23050_ (.A(\latched_rd[2] ),
    .B(\latched_rd[3] ),
    .C(_19366_),
    .X(_19560_));
 sky130_fd_sc_hd__nor2_1 _23051_ (.A(_19560_),
    .B(_19372_),
    .Y(_19561_));
 sky130_fd_sc_hd__buf_6 _23052_ (.A(_19561_),
    .X(_19562_));
 sky130_fd_sc_hd__clkbuf_4 _23053_ (.A(_19562_),
    .X(_19563_));
 sky130_fd_sc_hd__mux2_1 _23054_ (.A0(\cpuregs[16][31] ),
    .A1(\cpuregs_wrdata[31] ),
    .S(_19563_),
    .X(_03342_));
 sky130_fd_sc_hd__mux2_1 _23055_ (.A0(\cpuregs[16][30] ),
    .A1(\cpuregs_wrdata[30] ),
    .S(_19563_),
    .X(_03341_));
 sky130_fd_sc_hd__mux2_1 _23056_ (.A0(\cpuregs[16][29] ),
    .A1(\cpuregs_wrdata[29] ),
    .S(_19563_),
    .X(_03340_));
 sky130_fd_sc_hd__mux2_1 _23057_ (.A0(\cpuregs[16][28] ),
    .A1(\cpuregs_wrdata[28] ),
    .S(_19563_),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _23058_ (.A0(\cpuregs[16][27] ),
    .A1(\cpuregs_wrdata[27] ),
    .S(_19563_),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_1 _23059_ (.A0(\cpuregs[16][26] ),
    .A1(\cpuregs_wrdata[26] ),
    .S(_19563_),
    .X(_03337_));
 sky130_fd_sc_hd__buf_2 _23060_ (.A(_19562_),
    .X(_19564_));
 sky130_fd_sc_hd__mux2_1 _23061_ (.A0(\cpuregs[16][25] ),
    .A1(\cpuregs_wrdata[25] ),
    .S(_19564_),
    .X(_03336_));
 sky130_fd_sc_hd__mux2_1 _23062_ (.A0(\cpuregs[16][24] ),
    .A1(\cpuregs_wrdata[24] ),
    .S(_19564_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _23063_ (.A0(\cpuregs[16][23] ),
    .A1(\cpuregs_wrdata[23] ),
    .S(_19564_),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_1 _23064_ (.A0(\cpuregs[16][22] ),
    .A1(\cpuregs_wrdata[22] ),
    .S(_19564_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _23065_ (.A0(\cpuregs[16][21] ),
    .A1(\cpuregs_wrdata[21] ),
    .S(_19564_),
    .X(_03332_));
 sky130_fd_sc_hd__mux2_1 _23066_ (.A0(\cpuregs[16][20] ),
    .A1(\cpuregs_wrdata[20] ),
    .S(_19564_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_4 _23067_ (.A(_19562_),
    .X(_19565_));
 sky130_fd_sc_hd__mux2_1 _23068_ (.A0(\cpuregs[16][19] ),
    .A1(\cpuregs_wrdata[19] ),
    .S(_19565_),
    .X(_03330_));
 sky130_fd_sc_hd__mux2_1 _23069_ (.A0(\cpuregs[16][18] ),
    .A1(\cpuregs_wrdata[18] ),
    .S(_19565_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_1 _23070_ (.A0(\cpuregs[16][17] ),
    .A1(\cpuregs_wrdata[17] ),
    .S(_19565_),
    .X(_03328_));
 sky130_fd_sc_hd__mux2_1 _23071_ (.A0(\cpuregs[16][16] ),
    .A1(\cpuregs_wrdata[16] ),
    .S(_19565_),
    .X(_03327_));
 sky130_fd_sc_hd__mux2_1 _23072_ (.A0(\cpuregs[16][15] ),
    .A1(\cpuregs_wrdata[15] ),
    .S(_19565_),
    .X(_03326_));
 sky130_fd_sc_hd__mux2_1 _23073_ (.A0(\cpuregs[16][14] ),
    .A1(\cpuregs_wrdata[14] ),
    .S(_19565_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_4 _23074_ (.A(_19562_),
    .X(_19566_));
 sky130_fd_sc_hd__mux2_1 _23075_ (.A0(\cpuregs[16][13] ),
    .A1(\cpuregs_wrdata[13] ),
    .S(_19566_),
    .X(_03324_));
 sky130_fd_sc_hd__mux2_1 _23076_ (.A0(\cpuregs[16][12] ),
    .A1(\cpuregs_wrdata[12] ),
    .S(_19566_),
    .X(_03323_));
 sky130_fd_sc_hd__mux2_1 _23077_ (.A0(\cpuregs[16][11] ),
    .A1(\cpuregs_wrdata[11] ),
    .S(_19566_),
    .X(_03322_));
 sky130_fd_sc_hd__mux2_1 _23078_ (.A0(\cpuregs[16][10] ),
    .A1(\cpuregs_wrdata[10] ),
    .S(_19566_),
    .X(_03321_));
 sky130_fd_sc_hd__mux2_1 _23079_ (.A0(\cpuregs[16][9] ),
    .A1(\cpuregs_wrdata[9] ),
    .S(_19566_),
    .X(_03320_));
 sky130_fd_sc_hd__mux2_1 _23080_ (.A0(\cpuregs[16][8] ),
    .A1(\cpuregs_wrdata[8] ),
    .S(_19566_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_4 _23081_ (.A(_19561_),
    .X(_19567_));
 sky130_fd_sc_hd__mux2_1 _23082_ (.A0(\cpuregs[16][7] ),
    .A1(\cpuregs_wrdata[7] ),
    .S(_19567_),
    .X(_03318_));
 sky130_fd_sc_hd__mux2_1 _23083_ (.A0(\cpuregs[16][6] ),
    .A1(\cpuregs_wrdata[6] ),
    .S(_19567_),
    .X(_03317_));
 sky130_fd_sc_hd__mux2_1 _23084_ (.A0(\cpuregs[16][5] ),
    .A1(\cpuregs_wrdata[5] ),
    .S(_19567_),
    .X(_03316_));
 sky130_fd_sc_hd__mux2_1 _23085_ (.A0(\cpuregs[16][4] ),
    .A1(\cpuregs_wrdata[4] ),
    .S(_19567_),
    .X(_03315_));
 sky130_fd_sc_hd__mux2_1 _23086_ (.A0(\cpuregs[16][3] ),
    .A1(\cpuregs_wrdata[3] ),
    .S(_19567_),
    .X(_03314_));
 sky130_fd_sc_hd__mux2_1 _23087_ (.A0(\cpuregs[16][2] ),
    .A1(\cpuregs_wrdata[2] ),
    .S(_19567_),
    .X(_03313_));
 sky130_fd_sc_hd__mux2_1 _23088_ (.A0(\cpuregs[16][1] ),
    .A1(\cpuregs_wrdata[1] ),
    .S(_19562_),
    .X(_03312_));
 sky130_fd_sc_hd__mux2_1 _23089_ (.A0(\cpuregs[16][0] ),
    .A1(\cpuregs_wrdata[0] ),
    .S(_19562_),
    .X(_03311_));
 sky130_fd_sc_hd__nand2_1 _23090_ (.A(_19415_),
    .B(_19464_),
    .Y(_19568_));
 sky130_fd_sc_hd__buf_6 _23091_ (.A(_19568_),
    .X(_19569_));
 sky130_fd_sc_hd__clkbuf_4 _23092_ (.A(_19569_),
    .X(_19570_));
 sky130_fd_sc_hd__mux2_1 _23093_ (.A0(_19499_),
    .A1(\cpuregs[17][31] ),
    .S(_19570_),
    .X(_03310_));
 sky130_fd_sc_hd__mux2_1 _23094_ (.A0(_19503_),
    .A1(\cpuregs[17][30] ),
    .S(_19570_),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_1 _23095_ (.A0(_19504_),
    .A1(\cpuregs[17][29] ),
    .S(_19570_),
    .X(_03308_));
 sky130_fd_sc_hd__mux2_1 _23096_ (.A0(_19505_),
    .A1(\cpuregs[17][28] ),
    .S(_19570_),
    .X(_03307_));
 sky130_fd_sc_hd__mux2_1 _23097_ (.A0(_19506_),
    .A1(\cpuregs[17][27] ),
    .S(_19570_),
    .X(_03306_));
 sky130_fd_sc_hd__mux2_1 _23098_ (.A0(_19507_),
    .A1(\cpuregs[17][26] ),
    .S(_19570_),
    .X(_03305_));
 sky130_fd_sc_hd__buf_2 _23099_ (.A(_19569_),
    .X(_19571_));
 sky130_fd_sc_hd__mux2_1 _23100_ (.A0(_19508_),
    .A1(\cpuregs[17][25] ),
    .S(_19571_),
    .X(_03304_));
 sky130_fd_sc_hd__mux2_1 _23101_ (.A0(_19510_),
    .A1(\cpuregs[17][24] ),
    .S(_19571_),
    .X(_03303_));
 sky130_fd_sc_hd__mux2_1 _23102_ (.A0(_19511_),
    .A1(\cpuregs[17][23] ),
    .S(_19571_),
    .X(_03302_));
 sky130_fd_sc_hd__mux2_1 _23103_ (.A0(_19512_),
    .A1(\cpuregs[17][22] ),
    .S(_19571_),
    .X(_03301_));
 sky130_fd_sc_hd__mux2_1 _23104_ (.A0(_19513_),
    .A1(\cpuregs[17][21] ),
    .S(_19571_),
    .X(_03300_));
 sky130_fd_sc_hd__mux2_1 _23105_ (.A0(_19514_),
    .A1(\cpuregs[17][20] ),
    .S(_19571_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_4 _23106_ (.A(_19569_),
    .X(_19572_));
 sky130_fd_sc_hd__mux2_1 _23107_ (.A0(_19515_),
    .A1(\cpuregs[17][19] ),
    .S(_19572_),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_1 _23108_ (.A0(_19517_),
    .A1(\cpuregs[17][18] ),
    .S(_19572_),
    .X(_03297_));
 sky130_fd_sc_hd__mux2_1 _23109_ (.A0(_19518_),
    .A1(\cpuregs[17][17] ),
    .S(_19572_),
    .X(_03296_));
 sky130_fd_sc_hd__mux2_1 _23110_ (.A0(_19519_),
    .A1(\cpuregs[17][16] ),
    .S(_19572_),
    .X(_03295_));
 sky130_fd_sc_hd__mux2_1 _23111_ (.A0(_19520_),
    .A1(\cpuregs[17][15] ),
    .S(_19572_),
    .X(_03294_));
 sky130_fd_sc_hd__mux2_1 _23112_ (.A0(_19521_),
    .A1(\cpuregs[17][14] ),
    .S(_19572_),
    .X(_03293_));
 sky130_fd_sc_hd__buf_2 _23113_ (.A(_19569_),
    .X(_19573_));
 sky130_fd_sc_hd__mux2_1 _23114_ (.A0(_19522_),
    .A1(\cpuregs[17][13] ),
    .S(_19573_),
    .X(_03292_));
 sky130_fd_sc_hd__mux2_1 _23115_ (.A0(_19524_),
    .A1(\cpuregs[17][12] ),
    .S(_19573_),
    .X(_03291_));
 sky130_fd_sc_hd__mux2_1 _23116_ (.A0(_19525_),
    .A1(\cpuregs[17][11] ),
    .S(_19573_),
    .X(_03290_));
 sky130_fd_sc_hd__mux2_1 _23117_ (.A0(_19526_),
    .A1(\cpuregs[17][10] ),
    .S(_19573_),
    .X(_03289_));
 sky130_fd_sc_hd__mux2_1 _23118_ (.A0(_19527_),
    .A1(\cpuregs[17][9] ),
    .S(_19573_),
    .X(_03288_));
 sky130_fd_sc_hd__mux2_1 _23119_ (.A0(_19528_),
    .A1(\cpuregs[17][8] ),
    .S(_19573_),
    .X(_03287_));
 sky130_fd_sc_hd__clkbuf_4 _23120_ (.A(_19568_),
    .X(_19574_));
 sky130_fd_sc_hd__mux2_1 _23121_ (.A0(_19529_),
    .A1(\cpuregs[17][7] ),
    .S(_19574_),
    .X(_03286_));
 sky130_fd_sc_hd__mux2_1 _23122_ (.A0(_19531_),
    .A1(\cpuregs[17][6] ),
    .S(_19574_),
    .X(_03285_));
 sky130_fd_sc_hd__mux2_1 _23123_ (.A0(_19532_),
    .A1(\cpuregs[17][5] ),
    .S(_19574_),
    .X(_03284_));
 sky130_fd_sc_hd__mux2_1 _23124_ (.A0(_19533_),
    .A1(\cpuregs[17][4] ),
    .S(_19574_),
    .X(_03283_));
 sky130_fd_sc_hd__mux2_1 _23125_ (.A0(_19534_),
    .A1(\cpuregs[17][3] ),
    .S(_19574_),
    .X(_03282_));
 sky130_fd_sc_hd__mux2_1 _23126_ (.A0(_19535_),
    .A1(\cpuregs[17][2] ),
    .S(_19574_),
    .X(_03281_));
 sky130_fd_sc_hd__mux2_1 _23127_ (.A0(_19536_),
    .A1(\cpuregs[17][1] ),
    .S(_19569_),
    .X(_03280_));
 sky130_fd_sc_hd__mux2_1 _23128_ (.A0(_19537_),
    .A1(\cpuregs[17][0] ),
    .S(_19569_),
    .X(_03279_));
 sky130_fd_sc_hd__buf_4 _23129_ (.A(\pcpi_mul.rs2[31] ),
    .X(_19575_));
 sky130_fd_sc_hd__buf_6 _23130_ (.A(_19575_),
    .X(_19576_));
 sky130_fd_sc_hd__clkbuf_2 _23131_ (.A(_19576_),
    .X(_19577_));
 sky130_fd_sc_hd__clkbuf_2 _23132_ (.A(_19577_),
    .X(_19578_));
 sky130_fd_sc_hd__mux2_1 _23133_ (.A0(_19578_),
    .A1(_18471_),
    .S(_03728_),
    .X(_03278_));
 sky130_fd_sc_hd__clkbuf_2 _23134_ (.A(\pcpi_mul.rs2[30] ),
    .X(_19579_));
 sky130_fd_sc_hd__clkbuf_4 _23135_ (.A(net498),
    .X(_19580_));
 sky130_fd_sc_hd__buf_4 _23136_ (.A(_19580_),
    .X(_19581_));
 sky130_fd_sc_hd__mux2_1 _23137_ (.A0(_19581_),
    .A1(_19428_),
    .S(_03728_),
    .X(_03277_));
 sky130_fd_sc_hd__buf_4 _23138_ (.A(\pcpi_mul.rs2[29] ),
    .X(_19582_));
 sky130_fd_sc_hd__buf_6 _23139_ (.A(_19582_),
    .X(_19583_));
 sky130_fd_sc_hd__buf_2 _23140_ (.A(_19583_),
    .X(_19584_));
 sky130_fd_sc_hd__clkbuf_2 _23141_ (.A(_19584_),
    .X(_19585_));
 sky130_fd_sc_hd__mux2_1 _23142_ (.A0(_19585_),
    .A1(net359),
    .S(_03728_),
    .X(_03276_));
 sky130_fd_sc_hd__buf_4 _23143_ (.A(\pcpi_mul.rs2[28] ),
    .X(_19586_));
 sky130_fd_sc_hd__buf_6 _23144_ (.A(_19586_),
    .X(_19587_));
 sky130_fd_sc_hd__buf_4 _23145_ (.A(_19587_),
    .X(_19588_));
 sky130_fd_sc_hd__buf_2 _23146_ (.A(_19588_),
    .X(_19589_));
 sky130_fd_sc_hd__clkbuf_4 _23147_ (.A(_18464_),
    .X(_19590_));
 sky130_fd_sc_hd__mux2_1 _23148_ (.A0(_19589_),
    .A1(net358),
    .S(_19590_),
    .X(_03275_));
 sky130_fd_sc_hd__buf_4 _23149_ (.A(\pcpi_mul.rs2[27] ),
    .X(_19591_));
 sky130_fd_sc_hd__buf_6 _23150_ (.A(_19591_),
    .X(_19592_));
 sky130_fd_sc_hd__buf_6 _23151_ (.A(_19592_),
    .X(_19593_));
 sky130_fd_sc_hd__buf_2 _23152_ (.A(_19593_),
    .X(_19594_));
 sky130_fd_sc_hd__mux2_1 _23153_ (.A0(_19594_),
    .A1(_19429_),
    .S(_19590_),
    .X(_03274_));
 sky130_fd_sc_hd__clkbuf_4 _23154_ (.A(\pcpi_mul.rs2[26] ),
    .X(_19595_));
 sky130_fd_sc_hd__buf_4 _23155_ (.A(_19595_),
    .X(_19596_));
 sky130_fd_sc_hd__buf_4 _23156_ (.A(_19596_),
    .X(_19597_));
 sky130_fd_sc_hd__clkbuf_4 _23157_ (.A(_19597_),
    .X(_19598_));
 sky130_fd_sc_hd__mux2_1 _23158_ (.A0(_19598_),
    .A1(net356),
    .S(_19590_),
    .X(_03273_));
 sky130_fd_sc_hd__clkbuf_4 _23159_ (.A(\pcpi_mul.rs2[25] ),
    .X(_19599_));
 sky130_fd_sc_hd__buf_6 _23160_ (.A(_19599_),
    .X(_19600_));
 sky130_fd_sc_hd__clkbuf_4 _23161_ (.A(_19600_),
    .X(_19601_));
 sky130_fd_sc_hd__mux2_1 _23162_ (.A0(_19601_),
    .A1(net355),
    .S(_19590_),
    .X(_03272_));
 sky130_fd_sc_hd__buf_6 _23163_ (.A(\pcpi_mul.rs2[24] ),
    .X(_19602_));
 sky130_fd_sc_hd__buf_8 _23164_ (.A(_19602_),
    .X(_19603_));
 sky130_fd_sc_hd__buf_4 _23165_ (.A(_19603_),
    .X(_19604_));
 sky130_fd_sc_hd__clkbuf_4 _23166_ (.A(_19604_),
    .X(_19605_));
 sky130_fd_sc_hd__mux2_1 _23167_ (.A0(_19605_),
    .A1(net354),
    .S(_19590_),
    .X(_03271_));
 sky130_fd_sc_hd__buf_2 _23168_ (.A(\pcpi_mul.rs2[23] ),
    .X(_19606_));
 sky130_fd_sc_hd__buf_4 _23169_ (.A(_19606_),
    .X(_19607_));
 sky130_fd_sc_hd__buf_6 _23170_ (.A(_19607_),
    .X(_19608_));
 sky130_fd_sc_hd__buf_4 _23171_ (.A(_19608_),
    .X(_19609_));
 sky130_fd_sc_hd__mux2_1 _23172_ (.A0(_19609_),
    .A1(_19431_),
    .S(_19590_),
    .X(_03270_));
 sky130_fd_sc_hd__clkbuf_4 _23173_ (.A(\pcpi_mul.rs2[22] ),
    .X(_19610_));
 sky130_fd_sc_hd__buf_6 _23174_ (.A(_19610_),
    .X(_19611_));
 sky130_fd_sc_hd__buf_4 _23175_ (.A(_19611_),
    .X(_19612_));
 sky130_fd_sc_hd__buf_4 _23176_ (.A(_19612_),
    .X(_19613_));
 sky130_fd_sc_hd__buf_2 _23177_ (.A(_18464_),
    .X(_19614_));
 sky130_fd_sc_hd__mux2_1 _23178_ (.A0(_19613_),
    .A1(_19432_),
    .S(_19614_),
    .X(_03269_));
 sky130_fd_sc_hd__clkbuf_4 _23179_ (.A(\pcpi_mul.rs2[21] ),
    .X(_19615_));
 sky130_fd_sc_hd__buf_4 _23180_ (.A(_19615_),
    .X(_19616_));
 sky130_fd_sc_hd__clkbuf_8 _23181_ (.A(_19616_),
    .X(_19617_));
 sky130_fd_sc_hd__buf_2 _23182_ (.A(_19617_),
    .X(_19618_));
 sky130_fd_sc_hd__buf_4 _23183_ (.A(_19618_),
    .X(_19619_));
 sky130_fd_sc_hd__mux2_1 _23184_ (.A0(_19619_),
    .A1(_19433_),
    .S(_19614_),
    .X(_03268_));
 sky130_fd_sc_hd__buf_2 _23185_ (.A(\pcpi_mul.rs2[20] ),
    .X(_19620_));
 sky130_fd_sc_hd__buf_4 _23186_ (.A(_19620_),
    .X(_19621_));
 sky130_fd_sc_hd__buf_6 _23187_ (.A(_19621_),
    .X(_19622_));
 sky130_fd_sc_hd__clkbuf_4 _23188_ (.A(_19622_),
    .X(_19623_));
 sky130_fd_sc_hd__mux2_1 _23189_ (.A0(_19623_),
    .A1(net350),
    .S(_19614_),
    .X(_03267_));
 sky130_fd_sc_hd__buf_2 _23190_ (.A(\pcpi_mul.rs2[19] ),
    .X(_19624_));
 sky130_fd_sc_hd__clkbuf_8 _23191_ (.A(_19624_),
    .X(_19625_));
 sky130_fd_sc_hd__buf_6 _23192_ (.A(_19625_),
    .X(_19626_));
 sky130_fd_sc_hd__mux2_1 _23193_ (.A0(_19626_),
    .A1(net348),
    .S(_19614_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_6 _23194_ (.A(\pcpi_mul.rs2[18] ),
    .X(_19627_));
 sky130_fd_sc_hd__buf_4 _23195_ (.A(_19627_),
    .X(_19628_));
 sky130_fd_sc_hd__buf_4 _23196_ (.A(_19628_),
    .X(_19629_));
 sky130_fd_sc_hd__mux2_1 _23197_ (.A0(_19629_),
    .A1(_19435_),
    .S(_19614_),
    .X(_03265_));
 sky130_fd_sc_hd__clkbuf_2 _23198_ (.A(\pcpi_mul.rs2[17] ),
    .X(_19630_));
 sky130_fd_sc_hd__buf_6 _23199_ (.A(_19630_),
    .X(_19631_));
 sky130_fd_sc_hd__buf_4 _23200_ (.A(_19631_),
    .X(_19632_));
 sky130_fd_sc_hd__buf_6 _23201_ (.A(_19632_),
    .X(_19633_));
 sky130_fd_sc_hd__mux2_1 _23202_ (.A0(_19633_),
    .A1(net346),
    .S(_19614_),
    .X(_03264_));
 sky130_fd_sc_hd__buf_4 _23203_ (.A(\pcpi_mul.rs2[16] ),
    .X(_19634_));
 sky130_fd_sc_hd__buf_8 _23204_ (.A(_19634_),
    .X(_19635_));
 sky130_fd_sc_hd__buf_4 _23205_ (.A(_19635_),
    .X(_19636_));
 sky130_fd_sc_hd__clkbuf_8 _23206_ (.A(_19636_),
    .X(_19637_));
 sky130_fd_sc_hd__clkbuf_4 _23207_ (.A(_18463_),
    .X(_19638_));
 sky130_fd_sc_hd__buf_2 _23208_ (.A(_19638_),
    .X(_19639_));
 sky130_fd_sc_hd__mux2_1 _23209_ (.A0(_19637_),
    .A1(_19436_),
    .S(_19639_),
    .X(_03263_));
 sky130_fd_sc_hd__buf_6 _23210_ (.A(\pcpi_mul.rs2[15] ),
    .X(_19640_));
 sky130_fd_sc_hd__buf_4 _23211_ (.A(_19640_),
    .X(_19641_));
 sky130_fd_sc_hd__clkbuf_4 _23212_ (.A(_19641_),
    .X(_19642_));
 sky130_fd_sc_hd__mux2_1 _23213_ (.A0(net458),
    .A1(_19437_),
    .S(_19639_),
    .X(_03262_));
 sky130_fd_sc_hd__buf_4 _23214_ (.A(\pcpi_mul.rs2[14] ),
    .X(_19643_));
 sky130_fd_sc_hd__buf_6 _23215_ (.A(_19643_),
    .X(_19644_));
 sky130_fd_sc_hd__buf_4 _23216_ (.A(_19644_),
    .X(_19645_));
 sky130_fd_sc_hd__mux2_1 _23217_ (.A0(_19645_),
    .A1(_19438_),
    .S(_19639_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_4 _23218_ (.A(\pcpi_mul.rs2[13] ),
    .X(_19646_));
 sky130_fd_sc_hd__buf_6 _23219_ (.A(_19646_),
    .X(_19647_));
 sky130_fd_sc_hd__buf_6 _23220_ (.A(_19647_),
    .X(_19648_));
 sky130_fd_sc_hd__mux2_1 _23221_ (.A0(_19648_),
    .A1(_19440_),
    .S(_19639_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_4 _23222_ (.A(\pcpi_mul.rs2[12] ),
    .X(_19649_));
 sky130_fd_sc_hd__buf_2 _23223_ (.A(_19649_),
    .X(_19650_));
 sky130_fd_sc_hd__mux2_1 _23224_ (.A0(net478),
    .A1(_19441_),
    .S(_19639_),
    .X(_03259_));
 sky130_fd_sc_hd__clkbuf_4 _23225_ (.A(\pcpi_mul.rs2[11] ),
    .X(_19651_));
 sky130_fd_sc_hd__buf_1 _23226_ (.A(_19651_),
    .X(_19652_));
 sky130_fd_sc_hd__buf_8 _23227_ (.A(net477),
    .X(_19653_));
 sky130_fd_sc_hd__mux2_1 _23228_ (.A0(_19653_),
    .A1(_19442_),
    .S(_19639_),
    .X(_03258_));
 sky130_fd_sc_hd__clkbuf_4 _23229_ (.A(\pcpi_mul.rs2[10] ),
    .X(_19654_));
 sky130_fd_sc_hd__buf_6 _23230_ (.A(_19654_),
    .X(_19655_));
 sky130_fd_sc_hd__clkbuf_4 _23231_ (.A(_19655_),
    .X(_19656_));
 sky130_fd_sc_hd__buf_2 _23232_ (.A(_19638_),
    .X(_19657_));
 sky130_fd_sc_hd__mux2_1 _23233_ (.A0(net457),
    .A1(_19443_),
    .S(_19657_),
    .X(_03257_));
 sky130_fd_sc_hd__buf_6 _23234_ (.A(\pcpi_mul.rs2[9] ),
    .X(_19658_));
 sky130_fd_sc_hd__buf_8 _23235_ (.A(_19658_),
    .X(_19659_));
 sky130_fd_sc_hd__buf_1 _23236_ (.A(_19659_),
    .X(_19660_));
 sky130_fd_sc_hd__mux2_1 _23237_ (.A0(net456),
    .A1(_19444_),
    .S(_19657_),
    .X(_03256_));
 sky130_fd_sc_hd__buf_4 _23238_ (.A(\pcpi_mul.rs2[8] ),
    .X(_19661_));
 sky130_fd_sc_hd__buf_4 _23239_ (.A(_19661_),
    .X(_19662_));
 sky130_fd_sc_hd__buf_6 _23240_ (.A(_19662_),
    .X(_19663_));
 sky130_fd_sc_hd__mux2_1 _23241_ (.A0(_19663_),
    .A1(_19445_),
    .S(_19657_),
    .X(_03255_));
 sky130_fd_sc_hd__clkbuf_8 _23242_ (.A(\pcpi_mul.rs2[7] ),
    .X(_19664_));
 sky130_fd_sc_hd__buf_6 _23243_ (.A(_19664_),
    .X(_19665_));
 sky130_fd_sc_hd__buf_4 _23244_ (.A(_19665_),
    .X(_19666_));
 sky130_fd_sc_hd__mux2_1 _23245_ (.A0(_19666_),
    .A1(net499),
    .S(_19657_),
    .X(_03254_));
 sky130_fd_sc_hd__buf_6 _23246_ (.A(\pcpi_mul.rs2[6] ),
    .X(_19667_));
 sky130_fd_sc_hd__clkbuf_8 _23247_ (.A(_19667_),
    .X(_19668_));
 sky130_fd_sc_hd__mux2_1 _23248_ (.A0(_19668_),
    .A1(_19448_),
    .S(_19657_),
    .X(_03253_));
 sky130_fd_sc_hd__buf_6 _23249_ (.A(\pcpi_mul.rs2[5] ),
    .X(_19669_));
 sky130_fd_sc_hd__buf_6 _23250_ (.A(_19669_),
    .X(_19670_));
 sky130_fd_sc_hd__buf_2 _23251_ (.A(_19670_),
    .X(_19671_));
 sky130_fd_sc_hd__mux2_1 _23252_ (.A0(net455),
    .A1(_19449_),
    .S(_19657_),
    .X(_03252_));
 sky130_fd_sc_hd__buf_4 _23253_ (.A(\pcpi_mul.rs2[4] ),
    .X(_19672_));
 sky130_fd_sc_hd__buf_6 _23254_ (.A(_19672_),
    .X(_19673_));
 sky130_fd_sc_hd__buf_6 _23255_ (.A(_19673_),
    .X(_19674_));
 sky130_fd_sc_hd__buf_6 _23256_ (.A(_19638_),
    .X(_19675_));
 sky130_fd_sc_hd__mux2_1 _23257_ (.A0(_19674_),
    .A1(_19450_),
    .S(_19675_),
    .X(_03251_));
 sky130_fd_sc_hd__clkbuf_4 _23258_ (.A(\pcpi_mul.rs2[3] ),
    .X(_19676_));
 sky130_fd_sc_hd__buf_6 _23259_ (.A(_19676_),
    .X(_19677_));
 sky130_fd_sc_hd__mux2_1 _23260_ (.A0(_19677_),
    .A1(_19451_),
    .S(_19675_),
    .X(_03250_));
 sky130_fd_sc_hd__buf_4 _23261_ (.A(\pcpi_mul.rs2[2] ),
    .X(_19678_));
 sky130_fd_sc_hd__buf_6 _23262_ (.A(_19678_),
    .X(_19679_));
 sky130_fd_sc_hd__buf_4 _23263_ (.A(_19679_),
    .X(_19680_));
 sky130_fd_sc_hd__mux2_1 _23264_ (.A0(_19680_),
    .A1(_19452_),
    .S(_19675_),
    .X(_03249_));
 sky130_fd_sc_hd__buf_6 _23265_ (.A(\pcpi_mul.rs2[1] ),
    .X(_19681_));
 sky130_fd_sc_hd__clkbuf_4 _23266_ (.A(_19681_),
    .X(_19682_));
 sky130_fd_sc_hd__buf_6 _23267_ (.A(_19682_),
    .X(_19683_));
 sky130_fd_sc_hd__buf_4 _23268_ (.A(_19683_),
    .X(_19684_));
 sky130_fd_sc_hd__mux2_1 _23269_ (.A0(_19684_),
    .A1(_19453_),
    .S(_19675_),
    .X(_03248_));
 sky130_fd_sc_hd__buf_4 _23270_ (.A(\pcpi_mul.rs2[0] ),
    .X(_19685_));
 sky130_fd_sc_hd__buf_1 _23271_ (.A(_19685_),
    .X(_19686_));
 sky130_fd_sc_hd__buf_4 _23272_ (.A(net476),
    .X(_19687_));
 sky130_fd_sc_hd__mux2_1 _23273_ (.A0(_19687_),
    .A1(_19454_),
    .S(_19675_),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_1 _23274_ (.A0(net273),
    .A1(_02541_),
    .S(_18358_),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _23275_ (.A0(net272),
    .A1(_02540_),
    .S(_18358_),
    .X(_03245_));
 sky130_fd_sc_hd__mux2_1 _23276_ (.A0(net271),
    .A1(_02539_),
    .S(_18357_),
    .X(_03244_));
 sky130_fd_sc_hd__mux2_1 _23277_ (.A0(net270),
    .A1(_02538_),
    .S(_18357_),
    .X(_03243_));
 sky130_vsdinv _23278_ (.A(_00330_),
    .Y(_19688_));
 sky130_fd_sc_hd__and4_1 _23279_ (.A(_18365_),
    .B(_18369_),
    .C(_19688_),
    .D(_18371_),
    .X(_19689_));
 sky130_fd_sc_hd__clkbuf_2 _23280_ (.A(_18638_),
    .X(_19690_));
 sky130_fd_sc_hd__a32o_1 _23281_ (.A1(_19689_),
    .A2(_00329_),
    .A3(_00328_),
    .B1(is_alu_reg_reg),
    .B2(_19690_),
    .X(_03242_));
 sky130_vsdinv _23282_ (.A(_00329_),
    .Y(_19691_));
 sky130_fd_sc_hd__a32o_1 _23283_ (.A1(_19689_),
    .A2(_19691_),
    .A3(_00328_),
    .B1(is_alu_reg_imm),
    .B2(_19690_),
    .X(_03241_));
 sky130_fd_sc_hd__nand2_2 _23284_ (.A(_19415_),
    .B(_19491_),
    .Y(_19692_));
 sky130_fd_sc_hd__buf_8 _23285_ (.A(_19692_),
    .X(_19693_));
 sky130_fd_sc_hd__clkbuf_4 _23286_ (.A(_19693_),
    .X(_19694_));
 sky130_fd_sc_hd__mux2_1 _23287_ (.A0(_19499_),
    .A1(\cpuregs[13][31] ),
    .S(_19694_),
    .X(_03240_));
 sky130_fd_sc_hd__mux2_1 _23288_ (.A0(_19503_),
    .A1(\cpuregs[13][30] ),
    .S(_19694_),
    .X(_03239_));
 sky130_fd_sc_hd__mux2_1 _23289_ (.A0(_19504_),
    .A1(\cpuregs[13][29] ),
    .S(_19694_),
    .X(_03238_));
 sky130_fd_sc_hd__mux2_1 _23290_ (.A0(_19505_),
    .A1(\cpuregs[13][28] ),
    .S(_19694_),
    .X(_03237_));
 sky130_fd_sc_hd__mux2_1 _23291_ (.A0(_19506_),
    .A1(\cpuregs[13][27] ),
    .S(_19694_),
    .X(_03236_));
 sky130_fd_sc_hd__mux2_1 _23292_ (.A0(_19507_),
    .A1(\cpuregs[13][26] ),
    .S(_19694_),
    .X(_03235_));
 sky130_fd_sc_hd__buf_2 _23293_ (.A(_19693_),
    .X(_19695_));
 sky130_fd_sc_hd__mux2_1 _23294_ (.A0(_19508_),
    .A1(\cpuregs[13][25] ),
    .S(_19695_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _23295_ (.A0(_19510_),
    .A1(\cpuregs[13][24] ),
    .S(_19695_),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_1 _23296_ (.A0(_19511_),
    .A1(\cpuregs[13][23] ),
    .S(_19695_),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _23297_ (.A0(_19512_),
    .A1(\cpuregs[13][22] ),
    .S(_19695_),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_1 _23298_ (.A0(_19513_),
    .A1(\cpuregs[13][21] ),
    .S(_19695_),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _23299_ (.A0(_19514_),
    .A1(\cpuregs[13][20] ),
    .S(_19695_),
    .X(_03229_));
 sky130_fd_sc_hd__clkbuf_4 _23300_ (.A(_19693_),
    .X(_19696_));
 sky130_fd_sc_hd__mux2_1 _23301_ (.A0(_19515_),
    .A1(\cpuregs[13][19] ),
    .S(_19696_),
    .X(_03228_));
 sky130_fd_sc_hd__mux2_1 _23302_ (.A0(_19517_),
    .A1(\cpuregs[13][18] ),
    .S(_19696_),
    .X(_03227_));
 sky130_fd_sc_hd__mux2_1 _23303_ (.A0(_19518_),
    .A1(\cpuregs[13][17] ),
    .S(_19696_),
    .X(_03226_));
 sky130_fd_sc_hd__mux2_1 _23304_ (.A0(_19519_),
    .A1(\cpuregs[13][16] ),
    .S(_19696_),
    .X(_03225_));
 sky130_fd_sc_hd__mux2_1 _23305_ (.A0(_19520_),
    .A1(\cpuregs[13][15] ),
    .S(_19696_),
    .X(_03224_));
 sky130_fd_sc_hd__mux2_1 _23306_ (.A0(_19521_),
    .A1(\cpuregs[13][14] ),
    .S(_19696_),
    .X(_03223_));
 sky130_fd_sc_hd__buf_2 _23307_ (.A(_19693_),
    .X(_19697_));
 sky130_fd_sc_hd__mux2_1 _23308_ (.A0(_19522_),
    .A1(\cpuregs[13][13] ),
    .S(_19697_),
    .X(_03222_));
 sky130_fd_sc_hd__mux2_1 _23309_ (.A0(_19524_),
    .A1(\cpuregs[13][12] ),
    .S(_19697_),
    .X(_03221_));
 sky130_fd_sc_hd__mux2_1 _23310_ (.A0(_19525_),
    .A1(\cpuregs[13][11] ),
    .S(_19697_),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_1 _23311_ (.A0(_19526_),
    .A1(\cpuregs[13][10] ),
    .S(_19697_),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_1 _23312_ (.A0(_19527_),
    .A1(\cpuregs[13][9] ),
    .S(_19697_),
    .X(_03218_));
 sky130_fd_sc_hd__mux2_1 _23313_ (.A0(_19528_),
    .A1(\cpuregs[13][8] ),
    .S(_19697_),
    .X(_03217_));
 sky130_fd_sc_hd__clkbuf_4 _23314_ (.A(_19692_),
    .X(_19698_));
 sky130_fd_sc_hd__mux2_1 _23315_ (.A0(_19529_),
    .A1(\cpuregs[13][7] ),
    .S(_19698_),
    .X(_03216_));
 sky130_fd_sc_hd__mux2_1 _23316_ (.A0(_19531_),
    .A1(\cpuregs[13][6] ),
    .S(_19698_),
    .X(_03215_));
 sky130_fd_sc_hd__mux2_1 _23317_ (.A0(_19532_),
    .A1(\cpuregs[13][5] ),
    .S(_19698_),
    .X(_03214_));
 sky130_fd_sc_hd__mux2_1 _23318_ (.A0(_19533_),
    .A1(\cpuregs[13][4] ),
    .S(_19698_),
    .X(_03213_));
 sky130_fd_sc_hd__mux2_1 _23319_ (.A0(_19534_),
    .A1(\cpuregs[13][3] ),
    .S(_19698_),
    .X(_03212_));
 sky130_fd_sc_hd__mux2_1 _23320_ (.A0(_19535_),
    .A1(\cpuregs[13][2] ),
    .S(_19698_),
    .X(_03211_));
 sky130_fd_sc_hd__mux2_1 _23321_ (.A0(_19536_),
    .A1(\cpuregs[13][1] ),
    .S(_19693_),
    .X(_03210_));
 sky130_fd_sc_hd__mux2_1 _23322_ (.A0(_19537_),
    .A1(\cpuregs[13][0] ),
    .S(_19693_),
    .X(_03209_));
 sky130_fd_sc_hd__a32o_1 _23323_ (.A1(_19689_),
    .A2(_00329_),
    .A3(_18636_),
    .B1(is_sb_sh_sw),
    .B2(_19690_),
    .X(_03208_));
 sky130_fd_sc_hd__buf_2 _23324_ (.A(_18728_),
    .X(_19699_));
 sky130_fd_sc_hd__buf_2 _23325_ (.A(_18645_),
    .X(_19700_));
 sky130_fd_sc_hd__clkbuf_4 _23326_ (.A(_19700_),
    .X(_19701_));
 sky130_fd_sc_hd__inv_2 _23327_ (.A(instr_jalr),
    .Y(_02063_));
 sky130_fd_sc_hd__nand2_1 _23328_ (.A(_19701_),
    .B(_02063_),
    .Y(_19702_));
 sky130_vsdinv _23329_ (.A(_00335_),
    .Y(_19703_));
 sky130_fd_sc_hd__o21a_1 _23330_ (.A1(_19703_),
    .A2(_18693_),
    .B1(is_alu_reg_imm),
    .X(_19704_));
 sky130_fd_sc_hd__o22a_1 _23331_ (.A1(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .A2(_19699_),
    .B1(_19702_),
    .B2(_19704_),
    .X(_03207_));
 sky130_fd_sc_hd__o211a_1 _23332_ (.A1(_18659_),
    .A2(_18667_),
    .B1(_18660_),
    .C1(_18657_),
    .X(_19705_));
 sky130_fd_sc_hd__and3_1 _23333_ (.A(_18708_),
    .B(_18650_),
    .C(_18692_),
    .X(_19706_));
 sky130_fd_sc_hd__buf_4 _23334_ (.A(is_slli_srli_srai),
    .X(_19707_));
 sky130_fd_sc_hd__buf_2 _23335_ (.A(_18690_),
    .X(_19708_));
 sky130_fd_sc_hd__a32o_1 _23336_ (.A1(_19705_),
    .A2(_19706_),
    .A3(_18658_),
    .B1(_19707_),
    .B2(_19708_),
    .X(_03206_));
 sky130_fd_sc_hd__a32o_1 _23337_ (.A1(_19689_),
    .A2(_19691_),
    .A3(_18636_),
    .B1(is_lb_lh_lw_lbu_lhu),
    .B2(_19690_),
    .X(_03205_));
 sky130_fd_sc_hd__buf_4 _23338_ (.A(\decoded_imm_uj[20] ),
    .X(_19709_));
 sky130_fd_sc_hd__clkbuf_4 _23339_ (.A(_19709_),
    .X(_19710_));
 sky130_fd_sc_hd__buf_4 _23340_ (.A(_19710_),
    .X(_19711_));
 sky130_fd_sc_hd__mux2_4 _23341_ (.A0(_19711_),
    .A1(\mem_rdata_latched[31] ),
    .S(_18375_),
    .X(_03204_));
 sky130_fd_sc_hd__mux2_1 _23342_ (.A0(\decoded_imm_uj[19] ),
    .A1(\mem_rdata_latched[19] ),
    .S(_18375_),
    .X(_03203_));
 sky130_vsdinv _23343_ (.A(\decoded_imm_uj[18] ),
    .Y(_19712_));
 sky130_fd_sc_hd__o21ai_1 _23344_ (.A1(_19712_),
    .A2(_20895_),
    .B1(_18640_),
    .Y(_03202_));
 sky130_vsdinv _23345_ (.A(\decoded_imm_uj[17] ),
    .Y(_19713_));
 sky130_fd_sc_hd__o21ai_1 _23346_ (.A1(_19713_),
    .A2(_20895_),
    .B1(_18641_),
    .Y(_03201_));
 sky130_vsdinv _23347_ (.A(\decoded_imm_uj[16] ),
    .Y(_19714_));
 sky130_fd_sc_hd__o21ai_1 _23348_ (.A1(_19714_),
    .A2(_20895_),
    .B1(_18642_),
    .Y(_03200_));
 sky130_vsdinv _23349_ (.A(\decoded_imm_uj[15] ),
    .Y(_19715_));
 sky130_fd_sc_hd__o21ai_1 _23350_ (.A1(_19715_),
    .A2(_20895_),
    .B1(_18643_),
    .Y(_03199_));
 sky130_fd_sc_hd__clkbuf_4 _23351_ (.A(_18365_),
    .X(_19716_));
 sky130_fd_sc_hd__mux2_1 _23352_ (.A0(\decoded_imm_uj[14] ),
    .A1(\mem_rdata_latched[14] ),
    .S(_19716_),
    .X(_03198_));
 sky130_fd_sc_hd__mux2_1 _23353_ (.A0(\decoded_imm_uj[13] ),
    .A1(\mem_rdata_latched[13] ),
    .S(_19716_),
    .X(_03197_));
 sky130_fd_sc_hd__mux2_1 _23354_ (.A0(\decoded_imm_uj[12] ),
    .A1(\mem_rdata_latched[12] ),
    .S(_19716_),
    .X(_03196_));
 sky130_fd_sc_hd__mux2_1 _23355_ (.A0(\decoded_imm_uj[11] ),
    .A1(\mem_rdata_latched[20] ),
    .S(_19716_),
    .X(_03195_));
 sky130_fd_sc_hd__mux2_1 _23356_ (.A0(\decoded_imm_uj[10] ),
    .A1(\mem_rdata_latched[30] ),
    .S(_19716_),
    .X(_03194_));
 sky130_fd_sc_hd__mux2_1 _23357_ (.A0(\decoded_imm_uj[9] ),
    .A1(\mem_rdata_latched[29] ),
    .S(_19716_),
    .X(_03193_));
 sky130_fd_sc_hd__buf_2 _23358_ (.A(_18365_),
    .X(_19717_));
 sky130_fd_sc_hd__mux2_1 _23359_ (.A0(\decoded_imm_uj[8] ),
    .A1(\mem_rdata_latched[28] ),
    .S(_19717_),
    .X(_03192_));
 sky130_fd_sc_hd__and3_1 _23360_ (.A(_18361_),
    .B(_18346_),
    .C(\mem_rdata_latched[27] ),
    .X(_19718_));
 sky130_fd_sc_hd__a21o_1 _23361_ (.A1(_00337_),
    .A2(\decoded_imm_uj[7] ),
    .B1(_19718_),
    .X(_03191_));
 sky130_fd_sc_hd__mux2_1 _23362_ (.A0(\decoded_imm_uj[6] ),
    .A1(\mem_rdata_latched[26] ),
    .S(_19717_),
    .X(_03190_));
 sky130_fd_sc_hd__mux2_1 _23363_ (.A0(\decoded_imm_uj[5] ),
    .A1(\mem_rdata_latched[25] ),
    .S(_19717_),
    .X(_03189_));
 sky130_fd_sc_hd__mux2_1 _23364_ (.A0(\decoded_imm_uj[4] ),
    .A1(\mem_rdata_latched[24] ),
    .S(_19717_),
    .X(_03188_));
 sky130_fd_sc_hd__mux2_1 _23365_ (.A0(\decoded_imm_uj[3] ),
    .A1(\mem_rdata_latched[23] ),
    .S(_19717_),
    .X(_03187_));
 sky130_fd_sc_hd__mux2_1 _23366_ (.A0(\decoded_imm_uj[2] ),
    .A1(\mem_rdata_latched[22] ),
    .S(_19717_),
    .X(_03186_));
 sky130_fd_sc_hd__buf_2 _23367_ (.A(_18365_),
    .X(_19719_));
 sky130_fd_sc_hd__mux2_1 _23368_ (.A0(\decoded_imm_uj[1] ),
    .A1(\mem_rdata_latched[21] ),
    .S(_19719_),
    .X(_03185_));
 sky130_vsdinv _23369_ (.A(\mem_rdata_q[20] ),
    .Y(_19720_));
 sky130_vsdinv _23370_ (.A(is_alu_reg_imm),
    .Y(_19721_));
 sky130_fd_sc_hd__and3_1 _23371_ (.A(_19721_),
    .B(_18544_),
    .C(_02063_),
    .X(_19722_));
 sky130_fd_sc_hd__clkbuf_2 _23372_ (.A(_19722_),
    .X(_19723_));
 sky130_fd_sc_hd__a2bb2o_1 _23373_ (.A1_N(_19720_),
    .A2_N(_19723_),
    .B1(is_sb_sh_sw),
    .B2(\mem_rdata_q[7] ),
    .X(_19724_));
 sky130_fd_sc_hd__mux2_1 _23374_ (.A0(_19724_),
    .A1(\decoded_imm[0] ),
    .S(_18670_),
    .X(_03184_));
 sky130_fd_sc_hd__mux2_1 _23375_ (.A0(\decoded_rd[4] ),
    .A1(\mem_rdata_latched[11] ),
    .S(_19719_),
    .X(_03183_));
 sky130_fd_sc_hd__mux2_1 _23376_ (.A0(\decoded_rd[3] ),
    .A1(\mem_rdata_latched[10] ),
    .S(_19719_),
    .X(_03182_));
 sky130_fd_sc_hd__mux2_1 _23377_ (.A0(\decoded_rd[2] ),
    .A1(\mem_rdata_latched[9] ),
    .S(_19719_),
    .X(_03181_));
 sky130_fd_sc_hd__mux2_1 _23378_ (.A0(\decoded_rd[1] ),
    .A1(\mem_rdata_latched[8] ),
    .S(_19719_),
    .X(_03180_));
 sky130_fd_sc_hd__mux2_1 _23379_ (.A0(\decoded_rd[0] ),
    .A1(\mem_rdata_latched[7] ),
    .S(_19719_),
    .X(_03179_));
 sky130_fd_sc_hd__clkbuf_4 _23380_ (.A(instr_timer),
    .X(_19725_));
 sky130_fd_sc_hd__buf_2 _23381_ (.A(_18711_),
    .X(_19726_));
 sky130_fd_sc_hd__or3b_2 _23382_ (.A(\mem_rdata_q[4] ),
    .B(\mem_rdata_q[2] ),
    .C_N(\mem_rdata_q[3] ),
    .X(_19727_));
 sky130_fd_sc_hd__and2_1 _23383_ (.A(\mem_rdata_q[1] ),
    .B(\mem_rdata_q[0] ),
    .X(_19728_));
 sky130_fd_sc_hd__or4b_4 _23384_ (.A(\mem_rdata_q[6] ),
    .B(\mem_rdata_q[5] ),
    .C(_19727_),
    .D_N(_19728_),
    .X(_19729_));
 sky130_vsdinv _23385_ (.A(_19729_),
    .Y(_19730_));
 sky130_fd_sc_hd__and3_1 _23386_ (.A(_18661_),
    .B(\mem_rdata_q[25] ),
    .C(_18654_),
    .X(_19731_));
 sky130_fd_sc_hd__and3_1 _23387_ (.A(_19731_),
    .B(\mem_rdata_q[27] ),
    .C(_18728_),
    .X(_19732_));
 sky130_fd_sc_hd__a22o_1 _23388_ (.A1(_19725_),
    .A2(_19726_),
    .B1(_19730_),
    .B2(_19732_),
    .X(_03178_));
 sky130_fd_sc_hd__nor2_1 _23389_ (.A(_18368_),
    .B(_18372_),
    .Y(_19733_));
 sky130_fd_sc_hd__a22o_1 _23390_ (.A1(_19718_),
    .A2(_19733_),
    .B1(_19690_),
    .B2(instr_waitirq),
    .X(_03177_));
 sky130_fd_sc_hd__buf_2 _23391_ (.A(decoder_trigger),
    .X(_19734_));
 sky130_fd_sc_hd__and3_1 _23392_ (.A(_18655_),
    .B(_18707_),
    .C(_19734_),
    .X(_19735_));
 sky130_vsdinv _23393_ (.A(\mem_rdata_q[28] ),
    .Y(_19736_));
 sky130_fd_sc_hd__clkbuf_4 _23394_ (.A(\mem_rdata_q[26] ),
    .X(_19737_));
 sky130_fd_sc_hd__and4_1 _23395_ (.A(_18661_),
    .B(_19736_),
    .C(_19737_),
    .D(\mem_rdata_q[25] ),
    .X(_19738_));
 sky130_fd_sc_hd__clkbuf_4 _23396_ (.A(_18493_),
    .X(_19739_));
 sky130_fd_sc_hd__a32o_1 _23397_ (.A1(_19730_),
    .A2(_19735_),
    .A3(_19738_),
    .B1(_19739_),
    .B2(_19726_),
    .X(_03176_));
 sky130_fd_sc_hd__o21ai_1 _23398_ (.A1(_18339_),
    .A2(_18366_),
    .B1(_18380_),
    .Y(_03175_));
 sky130_fd_sc_hd__a32o_1 _23399_ (.A1(_19730_),
    .A2(_19731_),
    .A3(_19735_),
    .B1(instr_setq),
    .B2(_19726_),
    .X(_03174_));
 sky130_fd_sc_hd__clkbuf_2 _23400_ (.A(_18711_),
    .X(_19740_));
 sky130_fd_sc_hd__a22o_1 _23401_ (.A1(instr_getq),
    .A2(_19740_),
    .B1(_19730_),
    .B2(_18684_),
    .X(_03173_));
 sky130_fd_sc_hd__or4_1 _23402_ (.A(\mem_rdata_q[9] ),
    .B(\mem_rdata_q[8] ),
    .C(\mem_rdata_q[7] ),
    .D(_18703_),
    .X(_19741_));
 sky130_fd_sc_hd__nor2_1 _23403_ (.A(\mem_rdata_q[11] ),
    .B(\mem_rdata_q[10] ),
    .Y(_19742_));
 sky130_fd_sc_hd__nor2_1 _23404_ (.A(\mem_rdata_q[23] ),
    .B(\mem_rdata_q[22] ),
    .Y(_19743_));
 sky130_fd_sc_hd__nor2_1 _23405_ (.A(\mem_rdata_q[24] ),
    .B(\mem_rdata_q[21] ),
    .Y(_19744_));
 sky130_fd_sc_hd__and4b_1 _23406_ (.A_N(_19741_),
    .B(_19742_),
    .C(_19743_),
    .D(_19744_),
    .X(_19745_));
 sky130_fd_sc_hd__or2_1 _23407_ (.A(\mem_rdata_q[19] ),
    .B(\mem_rdata_q[18] ),
    .X(_19746_));
 sky130_fd_sc_hd__or4_4 _23408_ (.A(\mem_rdata_q[17] ),
    .B(\mem_rdata_q[16] ),
    .C(\mem_rdata_q[15] ),
    .D(_19746_),
    .X(_19747_));
 sky130_vsdinv _23409_ (.A(_19747_),
    .Y(_19748_));
 sky130_fd_sc_hd__or3b_2 _23410_ (.A(\mem_rdata_q[3] ),
    .B(\mem_rdata_q[2] ),
    .C_N(\mem_rdata_q[4] ),
    .X(_19749_));
 sky130_fd_sc_hd__and4b_1 _23411_ (.A_N(_19749_),
    .B(\mem_rdata_q[6] ),
    .C(\mem_rdata_q[5] ),
    .D(_19728_),
    .X(_19750_));
 sky130_fd_sc_hd__and3_1 _23412_ (.A(_19745_),
    .B(_19748_),
    .C(_19750_),
    .X(_19751_));
 sky130_fd_sc_hd__a22o_1 _23413_ (.A1(instr_ecall_ebreak),
    .A2(_19740_),
    .B1(_19751_),
    .B2(_18684_),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_2 _23414_ (.A(instr_rdinstrh),
    .X(_19752_));
 sky130_fd_sc_hd__and3_1 _23415_ (.A(_19748_),
    .B(_18698_),
    .C(_19743_),
    .X(_19753_));
 sky130_fd_sc_hd__and3_1 _23416_ (.A(_19720_),
    .B(_18707_),
    .C(_19734_),
    .X(_19754_));
 sky130_fd_sc_hd__and4_2 _23417_ (.A(_19753_),
    .B(\mem_rdata_q[21] ),
    .C(_19750_),
    .D(_19754_),
    .X(_19755_));
 sky130_fd_sc_hd__and3_1 _23418_ (.A(_18660_),
    .B(_19736_),
    .C(_18672_),
    .X(_19756_));
 sky130_fd_sc_hd__and3_1 _23419_ (.A(_19756_),
    .B(\mem_rdata_q[30] ),
    .C(_18656_),
    .X(_19757_));
 sky130_fd_sc_hd__nor2_1 _23420_ (.A(_19737_),
    .B(\mem_rdata_q[24] ),
    .Y(_19758_));
 sky130_fd_sc_hd__and3_1 _23421_ (.A(_19757_),
    .B(\mem_rdata_q[27] ),
    .C(_19758_),
    .X(_19759_));
 sky130_fd_sc_hd__a22o_1 _23422_ (.A1(_19752_),
    .A2(_19740_),
    .B1(_19755_),
    .B2(_19759_),
    .X(_03171_));
 sky130_fd_sc_hd__clkbuf_2 _23423_ (.A(instr_rdinstr),
    .X(_19760_));
 sky130_fd_sc_hd__clkbuf_4 _23424_ (.A(_19760_),
    .X(_19761_));
 sky130_fd_sc_hd__and3_1 _23425_ (.A(_19757_),
    .B(_18655_),
    .C(_19758_),
    .X(_19762_));
 sky130_fd_sc_hd__a22o_1 _23426_ (.A1(_19761_),
    .A2(_19740_),
    .B1(_19755_),
    .B2(_19762_),
    .X(_03170_));
 sky130_fd_sc_hd__clkbuf_4 _23427_ (.A(instr_rdcycleh),
    .X(_19763_));
 sky130_vsdinv _23428_ (.A(\mem_rdata_q[21] ),
    .Y(_19764_));
 sky130_fd_sc_hd__and3_1 _23429_ (.A(_19764_),
    .B(_18707_),
    .C(_19734_),
    .X(_19765_));
 sky130_fd_sc_hd__and3_1 _23430_ (.A(_19753_),
    .B(_19750_),
    .C(_19765_),
    .X(_19766_));
 sky130_fd_sc_hd__a22o_1 _23431_ (.A1(_19763_),
    .A2(_19740_),
    .B1(_19766_),
    .B2(_19759_),
    .X(_03169_));
 sky130_fd_sc_hd__a22o_1 _23432_ (.A1(instr_rdcycle),
    .A2(_19740_),
    .B1(_19766_),
    .B2(_19762_),
    .X(_03168_));
 sky130_fd_sc_hd__nor2_1 _23433_ (.A(_19721_),
    .B(_18679_),
    .Y(_19767_));
 sky130_fd_sc_hd__a22o_1 _23434_ (.A1(instr_srai),
    .A2(_18712_),
    .B1(_18677_),
    .B2(_19767_),
    .X(_03167_));
 sky130_fd_sc_hd__a22o_1 _23435_ (.A1(instr_srli),
    .A2(_18712_),
    .B1(_18684_),
    .B2(_19767_),
    .X(_03166_));
 sky130_fd_sc_hd__a32o_1 _23436_ (.A1(_18684_),
    .A2(is_alu_reg_imm),
    .A3(_18700_),
    .B1(instr_slli),
    .B2(_19726_),
    .X(_03165_));
 sky130_fd_sc_hd__and3_1 _23437_ (.A(_18707_),
    .B(is_sb_sh_sw),
    .C(_19734_),
    .X(_19768_));
 sky130_fd_sc_hd__a22o_1 _23438_ (.A1(instr_sw),
    .A2(_18712_),
    .B1(_18698_),
    .B2(_19768_),
    .X(_03164_));
 sky130_fd_sc_hd__a22o_1 _23439_ (.A1(_18700_),
    .A2(_19768_),
    .B1(_19708_),
    .B2(instr_sh),
    .X(_03163_));
 sky130_fd_sc_hd__a22o_1 _23440_ (.A1(_18702_),
    .A2(_19768_),
    .B1(instr_sb),
    .B2(_19726_),
    .X(_03162_));
 sky130_fd_sc_hd__and3_2 _23441_ (.A(_18707_),
    .B(is_lb_lh_lw_lbu_lhu),
    .C(_19734_),
    .X(_19769_));
 sky130_fd_sc_hd__a22o_1 _23442_ (.A1(_18678_),
    .A2(_19769_),
    .B1(_19708_),
    .B2(instr_lhu),
    .X(_03161_));
 sky130_fd_sc_hd__a22o_1 _23443_ (.A1(_18688_),
    .A2(_19769_),
    .B1(_19708_),
    .B2(instr_lbu),
    .X(_03160_));
 sky130_fd_sc_hd__a22o_1 _23444_ (.A1(instr_lw),
    .A2(_18712_),
    .B1(_18698_),
    .B2(_19769_),
    .X(_03159_));
 sky130_fd_sc_hd__a22o_1 _23445_ (.A1(_18700_),
    .A2(_19769_),
    .B1(_19708_),
    .B2(instr_lh),
    .X(_03158_));
 sky130_fd_sc_hd__a22o_1 _23446_ (.A1(_18702_),
    .A2(_19769_),
    .B1(instr_lb),
    .B2(_19726_),
    .X(_03157_));
 sky130_fd_sc_hd__nor3_4 _23447_ (.A(\mem_rdata_latched[14] ),
    .B(\mem_rdata_latched[13] ),
    .C(\mem_rdata_latched[12] ),
    .Y(_19770_));
 sky130_fd_sc_hd__and3_1 _23448_ (.A(_00325_),
    .B(_00324_),
    .C(_00326_),
    .X(_19771_));
 sky130_fd_sc_hd__and2_1 _23449_ (.A(_19771_),
    .B(_18369_),
    .X(_19772_));
 sky130_fd_sc_hd__nor2_1 _23450_ (.A(_02063_),
    .B(_18364_),
    .Y(_19773_));
 sky130_fd_sc_hd__a41o_1 _23451_ (.A1(_18366_),
    .A2(_18637_),
    .A3(_19770_),
    .A4(_19772_),
    .B1(_19773_),
    .X(_03156_));
 sky130_fd_sc_hd__nor2_1 _23452_ (.A(_00323_),
    .B(_18364_),
    .Y(_19774_));
 sky130_fd_sc_hd__a41o_1 _23453_ (.A1(_00327_),
    .A2(_18366_),
    .A3(_18637_),
    .A4(_19771_),
    .B1(_19774_),
    .X(_03155_));
 sky130_fd_sc_hd__and3_1 _23454_ (.A(_18364_),
    .B(_19688_),
    .C(_19772_),
    .X(_19775_));
 sky130_fd_sc_hd__a32o_1 _23455_ (.A1(_19775_),
    .A2(_19691_),
    .A3(_00328_),
    .B1(instr_auipc),
    .B2(_19690_),
    .X(_03154_));
 sky130_fd_sc_hd__buf_4 _23456_ (.A(instr_lui),
    .X(_19776_));
 sky130_fd_sc_hd__a32o_1 _23457_ (.A1(_19775_),
    .A2(_00329_),
    .A3(_00328_),
    .B1(_19776_),
    .B2(_18638_),
    .X(_03153_));
 sky130_fd_sc_hd__mux2_1 _23458_ (.A0(net298),
    .A1(_18672_),
    .S(_19701_),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_1 _23459_ (.A0(net297),
    .A1(\mem_rdata_q[30] ),
    .S(_19701_),
    .X(_03151_));
 sky130_fd_sc_hd__buf_2 _23460_ (.A(_18728_),
    .X(_19777_));
 sky130_fd_sc_hd__o21a_1 _23461_ (.A1(net295),
    .A2(_19777_),
    .B1(_18675_),
    .X(_03150_));
 sky130_fd_sc_hd__mux2_1 _23462_ (.A0(net294),
    .A1(\mem_rdata_q[28] ),
    .S(_19701_),
    .X(_03149_));
 sky130_fd_sc_hd__o21ba_1 _23463_ (.A1(net293),
    .A2(_19699_),
    .B1_N(_19735_),
    .X(_03148_));
 sky130_fd_sc_hd__mux2_1 _23464_ (.A0(net292),
    .A1(_19737_),
    .S(_19701_),
    .X(_03147_));
 sky130_fd_sc_hd__buf_2 _23465_ (.A(_19700_),
    .X(_19778_));
 sky130_fd_sc_hd__mux2_1 _23466_ (.A0(net291),
    .A1(\mem_rdata_q[25] ),
    .S(_19778_),
    .X(_03146_));
 sky130_fd_sc_hd__mux2_1 _23467_ (.A0(net290),
    .A1(\mem_rdata_q[24] ),
    .S(_19778_),
    .X(_03145_));
 sky130_fd_sc_hd__mux2_1 _23468_ (.A0(net289),
    .A1(\mem_rdata_q[23] ),
    .S(_19778_),
    .X(_03144_));
 sky130_fd_sc_hd__mux2_1 _23469_ (.A0(net288),
    .A1(\mem_rdata_q[22] ),
    .S(_19778_),
    .X(_03143_));
 sky130_fd_sc_hd__o21ba_1 _23470_ (.A1(net287),
    .A2(_19699_),
    .B1_N(_19765_),
    .X(_03142_));
 sky130_fd_sc_hd__o21ba_1 _23471_ (.A1(net286),
    .A2(_19699_),
    .B1_N(_19754_),
    .X(_03141_));
 sky130_fd_sc_hd__mux2_1 _23472_ (.A0(net284),
    .A1(\mem_rdata_q[19] ),
    .S(_19778_),
    .X(_03140_));
 sky130_fd_sc_hd__mux2_1 _23473_ (.A0(net283),
    .A1(\mem_rdata_q[18] ),
    .S(_19778_),
    .X(_03139_));
 sky130_fd_sc_hd__buf_6 _23474_ (.A(_19700_),
    .X(_19779_));
 sky130_fd_sc_hd__mux2_1 _23475_ (.A0(net282),
    .A1(\mem_rdata_q[17] ),
    .S(_19779_),
    .X(_03138_));
 sky130_fd_sc_hd__mux2_1 _23476_ (.A0(net281),
    .A1(\mem_rdata_q[16] ),
    .S(_19779_),
    .X(_03137_));
 sky130_fd_sc_hd__mux2_1 _23477_ (.A0(net280),
    .A1(\mem_rdata_q[15] ),
    .S(_19779_),
    .X(_03136_));
 sky130_fd_sc_hd__mux2_1 _23478_ (.A0(net279),
    .A1(_18667_),
    .S(_19779_),
    .X(_03135_));
 sky130_fd_sc_hd__mux2_1 _23479_ (.A0(net278),
    .A1(\mem_rdata_q[13] ),
    .S(_19779_),
    .X(_03134_));
 sky130_fd_sc_hd__mux2_1 _23480_ (.A0(net277),
    .A1(_18692_),
    .S(_19779_),
    .X(_03133_));
 sky130_fd_sc_hd__buf_2 _23481_ (.A(_19700_),
    .X(_19780_));
 sky130_fd_sc_hd__mux2_1 _23482_ (.A0(net276),
    .A1(\mem_rdata_q[11] ),
    .S(_19780_),
    .X(_03132_));
 sky130_fd_sc_hd__mux2_1 _23483_ (.A0(net275),
    .A1(\mem_rdata_q[10] ),
    .S(_19780_),
    .X(_03131_));
 sky130_fd_sc_hd__mux2_1 _23484_ (.A0(net305),
    .A1(\mem_rdata_q[9] ),
    .S(_19780_),
    .X(_03130_));
 sky130_fd_sc_hd__mux2_1 _23485_ (.A0(net304),
    .A1(\mem_rdata_q[8] ),
    .S(_19780_),
    .X(_03129_));
 sky130_fd_sc_hd__mux2_1 _23486_ (.A0(net303),
    .A1(\mem_rdata_q[7] ),
    .S(_19780_),
    .X(_03128_));
 sky130_fd_sc_hd__mux2_1 _23487_ (.A0(net302),
    .A1(\mem_rdata_q[6] ),
    .S(_19780_),
    .X(_03127_));
 sky130_fd_sc_hd__buf_2 _23488_ (.A(_19700_),
    .X(_19781_));
 sky130_fd_sc_hd__mux2_1 _23489_ (.A0(net301),
    .A1(\mem_rdata_q[5] ),
    .S(_19781_),
    .X(_03126_));
 sky130_fd_sc_hd__mux2_1 _23490_ (.A0(net300),
    .A1(\mem_rdata_q[4] ),
    .S(_19781_),
    .X(_03125_));
 sky130_fd_sc_hd__mux2_1 _23491_ (.A0(net299),
    .A1(\mem_rdata_q[3] ),
    .S(_19781_),
    .X(_03124_));
 sky130_fd_sc_hd__mux2_1 _23492_ (.A0(net296),
    .A1(\mem_rdata_q[2] ),
    .S(_19781_),
    .X(_03123_));
 sky130_fd_sc_hd__mux2_1 _23493_ (.A0(net285),
    .A1(\mem_rdata_q[1] ),
    .S(_19781_),
    .X(_03122_));
 sky130_fd_sc_hd__mux2_1 _23494_ (.A0(net274),
    .A1(\mem_rdata_q[0] ),
    .S(_19781_),
    .X(_03121_));
 sky130_vsdinv _23495_ (.A(\cpu_state[5] ),
    .Y(_19782_));
 sky130_fd_sc_hd__or3_1 _23496_ (.A(_00318_),
    .B(_00320_),
    .C(_18309_),
    .X(_19783_));
 sky130_fd_sc_hd__a31o_2 _23497_ (.A1(_18541_),
    .A2(_18328_),
    .A3(_19782_),
    .B1(_19783_),
    .X(_19784_));
 sky130_fd_sc_hd__buf_2 _23498_ (.A(_19784_),
    .X(_19785_));
 sky130_fd_sc_hd__buf_2 _23499_ (.A(_19785_),
    .X(_19786_));
 sky130_fd_sc_hd__mux2_1 _23500_ (.A0(_02499_),
    .A1(_18451_),
    .S(_19786_),
    .X(_03120_));
 sky130_fd_sc_hd__clkbuf_4 _23501_ (.A(net329),
    .X(_19787_));
 sky130_fd_sc_hd__mux2_1 _23502_ (.A0(_02498_),
    .A1(_19787_),
    .S(_19786_),
    .X(_03119_));
 sky130_fd_sc_hd__buf_6 _23503_ (.A(net327),
    .X(_19788_));
 sky130_fd_sc_hd__mux2_1 _23504_ (.A0(_02496_),
    .A1(_19788_),
    .S(_19786_),
    .X(_03118_));
 sky130_fd_sc_hd__mux2_1 _23505_ (.A0(_02495_),
    .A1(net326),
    .S(_19786_),
    .X(_03117_));
 sky130_fd_sc_hd__buf_4 _23506_ (.A(net325),
    .X(_19789_));
 sky130_fd_sc_hd__mux2_1 _23507_ (.A0(_02494_),
    .A1(_19789_),
    .S(_19786_),
    .X(_03116_));
 sky130_fd_sc_hd__mux2_1 _23508_ (.A0(_02493_),
    .A1(net324),
    .S(_19786_),
    .X(_03115_));
 sky130_fd_sc_hd__buf_4 _23509_ (.A(net323),
    .X(_19790_));
 sky130_fd_sc_hd__buf_2 _23510_ (.A(_19785_),
    .X(_19791_));
 sky130_fd_sc_hd__mux2_1 _23511_ (.A0(_02492_),
    .A1(_19790_),
    .S(_19791_),
    .X(_03114_));
 sky130_fd_sc_hd__buf_4 _23512_ (.A(net322),
    .X(_19792_));
 sky130_fd_sc_hd__mux2_1 _23513_ (.A0(_02491_),
    .A1(_19792_),
    .S(_19791_),
    .X(_03113_));
 sky130_fd_sc_hd__buf_4 _23514_ (.A(net321),
    .X(_19793_));
 sky130_fd_sc_hd__mux2_1 _23515_ (.A0(_02490_),
    .A1(_19793_),
    .S(_19791_),
    .X(_03112_));
 sky130_fd_sc_hd__buf_4 _23516_ (.A(net320),
    .X(_19794_));
 sky130_fd_sc_hd__mux2_1 _23517_ (.A0(_02489_),
    .A1(_19794_),
    .S(_19791_),
    .X(_03111_));
 sky130_fd_sc_hd__buf_6 _23518_ (.A(net319),
    .X(_19795_));
 sky130_fd_sc_hd__mux2_1 _23519_ (.A0(_02488_),
    .A1(_19795_),
    .S(_19791_),
    .X(_03110_));
 sky130_fd_sc_hd__buf_4 _23520_ (.A(net318),
    .X(_19796_));
 sky130_fd_sc_hd__mux2_1 _23521_ (.A0(_02487_),
    .A1(_19796_),
    .S(_19791_),
    .X(_03109_));
 sky130_fd_sc_hd__buf_4 _23522_ (.A(net316),
    .X(_19797_));
 sky130_fd_sc_hd__buf_2 _23523_ (.A(_19785_),
    .X(_19798_));
 sky130_fd_sc_hd__mux2_1 _23524_ (.A0(_02485_),
    .A1(_19797_),
    .S(_19798_),
    .X(_03108_));
 sky130_fd_sc_hd__buf_4 _23525_ (.A(net315),
    .X(_19799_));
 sky130_fd_sc_hd__mux2_1 _23526_ (.A0(_02484_),
    .A1(_19799_),
    .S(_19798_),
    .X(_03107_));
 sky130_fd_sc_hd__buf_4 _23527_ (.A(net314),
    .X(_19800_));
 sky130_fd_sc_hd__mux2_1 _23528_ (.A0(_02483_),
    .A1(_19800_),
    .S(_19798_),
    .X(_03106_));
 sky130_fd_sc_hd__buf_4 _23529_ (.A(net313),
    .X(_19801_));
 sky130_fd_sc_hd__mux2_1 _23530_ (.A0(_02482_),
    .A1(_19801_),
    .S(_19798_),
    .X(_03105_));
 sky130_fd_sc_hd__buf_4 _23531_ (.A(net312),
    .X(_19802_));
 sky130_fd_sc_hd__mux2_1 _23532_ (.A0(_02481_),
    .A1(_19802_),
    .S(_19798_),
    .X(_03104_));
 sky130_fd_sc_hd__buf_4 _23533_ (.A(net311),
    .X(_19803_));
 sky130_fd_sc_hd__mux2_1 _23534_ (.A0(_02480_),
    .A1(_19803_),
    .S(_19798_),
    .X(_03103_));
 sky130_fd_sc_hd__buf_4 _23535_ (.A(net310),
    .X(_19804_));
 sky130_fd_sc_hd__buf_2 _23536_ (.A(_19785_),
    .X(_19805_));
 sky130_fd_sc_hd__mux2_1 _23537_ (.A0(_02479_),
    .A1(_19804_),
    .S(_19805_),
    .X(_03102_));
 sky130_fd_sc_hd__buf_4 _23538_ (.A(net309),
    .X(_19806_));
 sky130_fd_sc_hd__mux2_1 _23539_ (.A0(_02478_),
    .A1(_19806_),
    .S(_19805_),
    .X(_03101_));
 sky130_fd_sc_hd__buf_4 _23540_ (.A(net308),
    .X(_19807_));
 sky130_fd_sc_hd__mux2_1 _23541_ (.A0(_02477_),
    .A1(_19807_),
    .S(_19805_),
    .X(_03100_));
 sky130_fd_sc_hd__buf_4 _23542_ (.A(net307),
    .X(_19808_));
 sky130_fd_sc_hd__mux2_1 _23543_ (.A0(_02476_),
    .A1(_19808_),
    .S(_19805_),
    .X(_03099_));
 sky130_fd_sc_hd__buf_4 _23544_ (.A(net337),
    .X(_19809_));
 sky130_fd_sc_hd__mux2_1 _23545_ (.A0(_02506_),
    .A1(_19809_),
    .S(_19805_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_4 _23546_ (.A(net336),
    .X(_19810_));
 sky130_fd_sc_hd__mux2_1 _23547_ (.A0(_02505_),
    .A1(_19810_),
    .S(_19805_),
    .X(_03097_));
 sky130_fd_sc_hd__buf_4 _23548_ (.A(net335),
    .X(_19811_));
 sky130_fd_sc_hd__clkbuf_4 _23549_ (.A(_19784_),
    .X(_19812_));
 sky130_fd_sc_hd__mux2_1 _23550_ (.A0(_02504_),
    .A1(_19811_),
    .S(_19812_),
    .X(_03096_));
 sky130_fd_sc_hd__buf_6 _23551_ (.A(net334),
    .X(_19813_));
 sky130_fd_sc_hd__mux2_1 _23552_ (.A0(_02503_),
    .A1(_19813_),
    .S(_19812_),
    .X(_03095_));
 sky130_fd_sc_hd__buf_4 _23553_ (.A(net333),
    .X(_19814_));
 sky130_fd_sc_hd__mux2_1 _23554_ (.A0(_02502_),
    .A1(_19814_),
    .S(_19812_),
    .X(_03094_));
 sky130_fd_sc_hd__buf_4 _23555_ (.A(net332),
    .X(_19815_));
 sky130_fd_sc_hd__mux2_1 _23556_ (.A0(_02501_),
    .A1(_19815_),
    .S(_19812_),
    .X(_03093_));
 sky130_fd_sc_hd__buf_6 _23557_ (.A(net331),
    .X(_19816_));
 sky130_fd_sc_hd__mux2_1 _23558_ (.A0(_02500_),
    .A1(_19816_),
    .S(_19812_),
    .X(_03092_));
 sky130_fd_sc_hd__buf_4 _23559_ (.A(net328),
    .X(_19817_));
 sky130_fd_sc_hd__mux2_1 _23560_ (.A0(_02497_),
    .A1(_19817_),
    .S(_19812_),
    .X(_03091_));
 sky130_fd_sc_hd__buf_6 _23561_ (.A(net317),
    .X(_19818_));
 sky130_fd_sc_hd__buf_6 _23562_ (.A(_19818_),
    .X(_19819_));
 sky130_fd_sc_hd__mux2_1 _23563_ (.A0(_02486_),
    .A1(_19819_),
    .S(_19785_),
    .X(_03090_));
 sky130_fd_sc_hd__buf_6 _23564_ (.A(net306),
    .X(_19820_));
 sky130_fd_sc_hd__mux2_1 _23565_ (.A0(_02475_),
    .A1(_19820_),
    .S(_19785_),
    .X(_03089_));
 sky130_fd_sc_hd__mux2_1 _23566_ (.A0(net158),
    .A1(net191),
    .S(net422),
    .X(_03088_));
 sky130_fd_sc_hd__mux2_1 _23567_ (.A0(net157),
    .A1(net190),
    .S(_18635_),
    .X(_03087_));
 sky130_fd_sc_hd__mux2_1 _23568_ (.A0(net155),
    .A1(net188),
    .S(net422),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_1 _23569_ (.A0(net154),
    .A1(net187),
    .S(net422),
    .X(_03085_));
 sky130_fd_sc_hd__mux2_1 _23570_ (.A0(net153),
    .A1(net186),
    .S(_18635_),
    .X(_03084_));
 sky130_fd_sc_hd__clkbuf_4 _23571_ (.A(_18634_),
    .X(_19821_));
 sky130_fd_sc_hd__mux2_1 _23572_ (.A0(net152),
    .A1(net185),
    .S(net417),
    .X(_03083_));
 sky130_fd_sc_hd__mux2_1 _23573_ (.A0(net151),
    .A1(net184),
    .S(net417),
    .X(_03082_));
 sky130_fd_sc_hd__mux2_1 _23574_ (.A0(net150),
    .A1(net183),
    .S(net417),
    .X(_03081_));
 sky130_fd_sc_hd__mux2_1 _23575_ (.A0(net149),
    .A1(net182),
    .S(net417),
    .X(_03080_));
 sky130_fd_sc_hd__mux2_1 _23576_ (.A0(net148),
    .A1(net181),
    .S(_19821_),
    .X(_03079_));
 sky130_fd_sc_hd__mux2_1 _23577_ (.A0(net147),
    .A1(net180),
    .S(net417),
    .X(_03078_));
 sky130_fd_sc_hd__buf_6 _23578_ (.A(_18634_),
    .X(_19822_));
 sky130_fd_sc_hd__mux2_1 _23579_ (.A0(net146),
    .A1(net179),
    .S(net416),
    .X(_03077_));
 sky130_fd_sc_hd__mux2_1 _23580_ (.A0(net144),
    .A1(net177),
    .S(net416),
    .X(_03076_));
 sky130_fd_sc_hd__mux2_1 _23581_ (.A0(net143),
    .A1(net176),
    .S(net416),
    .X(_03075_));
 sky130_fd_sc_hd__mux2_1 _23582_ (.A0(net142),
    .A1(net175),
    .S(_19822_),
    .X(_03074_));
 sky130_fd_sc_hd__mux2_1 _23583_ (.A0(net141),
    .A1(net174),
    .S(_19822_),
    .X(_03073_));
 sky130_fd_sc_hd__mux2_1 _23584_ (.A0(net140),
    .A1(net173),
    .S(net416),
    .X(_03072_));
 sky130_fd_sc_hd__buf_8 _23585_ (.A(_18634_),
    .X(_19823_));
 sky130_fd_sc_hd__mux2_1 _23586_ (.A0(net139),
    .A1(net172),
    .S(_19823_),
    .X(_03071_));
 sky130_fd_sc_hd__mux2_1 _23587_ (.A0(net138),
    .A1(net171),
    .S(net415),
    .X(_03070_));
 sky130_fd_sc_hd__mux2_1 _23588_ (.A0(net137),
    .A1(net170),
    .S(net415),
    .X(_03069_));
 sky130_fd_sc_hd__mux2_1 _23589_ (.A0(net136),
    .A1(net169),
    .S(net415),
    .X(_03068_));
 sky130_fd_sc_hd__mux2_1 _23590_ (.A0(net135),
    .A1(net168),
    .S(_19823_),
    .X(_03067_));
 sky130_fd_sc_hd__mux2_1 _23591_ (.A0(net165),
    .A1(net198),
    .S(_19823_),
    .X(_03066_));
 sky130_fd_sc_hd__buf_4 _23592_ (.A(_18634_),
    .X(_19824_));
 sky130_fd_sc_hd__mux2_1 _23593_ (.A0(net164),
    .A1(net197),
    .S(net414),
    .X(_03065_));
 sky130_fd_sc_hd__mux2_1 _23594_ (.A0(net163),
    .A1(net196),
    .S(net414),
    .X(_03064_));
 sky130_fd_sc_hd__mux2_1 _23595_ (.A0(net162),
    .A1(net195),
    .S(net414),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_1 _23596_ (.A0(net161),
    .A1(net194),
    .S(net414),
    .X(_03062_));
 sky130_fd_sc_hd__mux2_1 _23597_ (.A0(net160),
    .A1(net193),
    .S(net414),
    .X(_03061_));
 sky130_fd_sc_hd__mux2_1 _23598_ (.A0(net159),
    .A1(net192),
    .S(_19824_),
    .X(_03060_));
 sky130_fd_sc_hd__mux2_1 _23599_ (.A0(net156),
    .A1(net189),
    .S(_18634_),
    .X(_03059_));
 sky130_fd_sc_hd__buf_4 _23600_ (.A(\pcpi_mul.rs1[31] ),
    .X(_19825_));
 sky130_fd_sc_hd__buf_6 _23601_ (.A(_19825_),
    .X(_19826_));
 sky130_fd_sc_hd__buf_6 _23602_ (.A(_19826_),
    .X(_19827_));
 sky130_fd_sc_hd__clkbuf_2 _23603_ (.A(_19827_),
    .X(_19828_));
 sky130_fd_sc_hd__mux2_1 _23604_ (.A0(_19828_),
    .A1(_18451_),
    .S(_19675_),
    .X(_03058_));
 sky130_fd_sc_hd__buf_4 _23605_ (.A(\pcpi_mul.rs1[30] ),
    .X(_19829_));
 sky130_fd_sc_hd__buf_6 _23606_ (.A(_19829_),
    .X(_19830_));
 sky130_fd_sc_hd__clkbuf_4 _23607_ (.A(_19830_),
    .X(_19831_));
 sky130_fd_sc_hd__buf_2 _23608_ (.A(_19831_),
    .X(_19832_));
 sky130_fd_sc_hd__clkbuf_4 _23609_ (.A(_19638_),
    .X(_19833_));
 sky130_fd_sc_hd__mux2_1 _23610_ (.A0(_19832_),
    .A1(_19787_),
    .S(_19833_),
    .X(_03057_));
 sky130_fd_sc_hd__buf_4 _23611_ (.A(\pcpi_mul.rs1[29] ),
    .X(_19834_));
 sky130_fd_sc_hd__buf_6 _23612_ (.A(_19834_),
    .X(_19835_));
 sky130_fd_sc_hd__buf_2 _23613_ (.A(_19835_),
    .X(_19836_));
 sky130_fd_sc_hd__clkbuf_4 _23614_ (.A(_19836_),
    .X(_19837_));
 sky130_fd_sc_hd__mux2_1 _23615_ (.A0(_19837_),
    .A1(_19788_),
    .S(_19833_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_4 _23616_ (.A(\pcpi_mul.rs1[28] ),
    .X(_19838_));
 sky130_fd_sc_hd__buf_4 _23617_ (.A(_19838_),
    .X(_19839_));
 sky130_fd_sc_hd__buf_4 _23618_ (.A(_19839_),
    .X(_19840_));
 sky130_fd_sc_hd__clkbuf_4 _23619_ (.A(_19840_),
    .X(_19841_));
 sky130_fd_sc_hd__buf_2 _23620_ (.A(_19841_),
    .X(_19842_));
 sky130_fd_sc_hd__mux2_1 _23621_ (.A0(_19842_),
    .A1(net326),
    .S(_19833_),
    .X(_03055_));
 sky130_fd_sc_hd__buf_6 _23622_ (.A(\pcpi_mul.rs1[27] ),
    .X(_19843_));
 sky130_fd_sc_hd__clkbuf_4 _23623_ (.A(_19843_),
    .X(_19844_));
 sky130_fd_sc_hd__clkbuf_4 _23624_ (.A(_19844_),
    .X(_19845_));
 sky130_fd_sc_hd__clkbuf_4 _23625_ (.A(_19845_),
    .X(_19846_));
 sky130_fd_sc_hd__mux2_1 _23626_ (.A0(_19846_),
    .A1(_19789_),
    .S(_19833_),
    .X(_03054_));
 sky130_fd_sc_hd__buf_2 _23627_ (.A(\pcpi_mul.rs1[26] ),
    .X(_19847_));
 sky130_fd_sc_hd__buf_4 _23628_ (.A(_19847_),
    .X(_19848_));
 sky130_fd_sc_hd__buf_4 _23629_ (.A(_19848_),
    .X(_19849_));
 sky130_fd_sc_hd__buf_4 _23630_ (.A(_19849_),
    .X(_19850_));
 sky130_fd_sc_hd__mux2_1 _23631_ (.A0(_19850_),
    .A1(net324),
    .S(_19833_),
    .X(_03053_));
 sky130_fd_sc_hd__buf_4 _23632_ (.A(\pcpi_mul.rs1[25] ),
    .X(_19851_));
 sky130_fd_sc_hd__clkbuf_2 _23633_ (.A(_19851_),
    .X(_19852_));
 sky130_fd_sc_hd__buf_4 _23634_ (.A(_19852_),
    .X(_19853_));
 sky130_fd_sc_hd__mux2_1 _23635_ (.A0(_19853_),
    .A1(_19790_),
    .S(_19833_),
    .X(_03052_));
 sky130_fd_sc_hd__buf_4 _23636_ (.A(\pcpi_mul.rs1[24] ),
    .X(_19854_));
 sky130_fd_sc_hd__buf_4 _23637_ (.A(_19854_),
    .X(_19855_));
 sky130_fd_sc_hd__buf_4 _23638_ (.A(_19855_),
    .X(_19856_));
 sky130_fd_sc_hd__clkbuf_4 _23639_ (.A(_19638_),
    .X(_19857_));
 sky130_fd_sc_hd__mux2_1 _23640_ (.A0(_19856_),
    .A1(_19792_),
    .S(_19857_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_4 _23641_ (.A(\pcpi_mul.rs1[23] ),
    .X(_19858_));
 sky130_fd_sc_hd__buf_6 _23642_ (.A(_19858_),
    .X(_19859_));
 sky130_fd_sc_hd__clkbuf_4 _23643_ (.A(_19859_),
    .X(_19860_));
 sky130_fd_sc_hd__mux2_1 _23644_ (.A0(_19860_),
    .A1(_19793_),
    .S(_19857_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_4 _23645_ (.A(\pcpi_mul.rs1[22] ),
    .X(_19861_));
 sky130_fd_sc_hd__buf_4 _23646_ (.A(_19861_),
    .X(_19862_));
 sky130_fd_sc_hd__buf_6 _23647_ (.A(_19862_),
    .X(_19863_));
 sky130_fd_sc_hd__buf_4 _23648_ (.A(_19863_),
    .X(_19864_));
 sky130_fd_sc_hd__mux2_1 _23649_ (.A0(_19864_),
    .A1(_19794_),
    .S(_19857_),
    .X(_03049_));
 sky130_fd_sc_hd__buf_6 _23650_ (.A(\pcpi_mul.rs1[21] ),
    .X(_19865_));
 sky130_fd_sc_hd__buf_4 _23651_ (.A(_19865_),
    .X(_19866_));
 sky130_fd_sc_hd__buf_4 _23652_ (.A(_19866_),
    .X(_19867_));
 sky130_fd_sc_hd__mux2_1 _23653_ (.A0(_19867_),
    .A1(_19795_),
    .S(_19857_),
    .X(_03048_));
 sky130_fd_sc_hd__buf_6 _23654_ (.A(\pcpi_mul.rs1[20] ),
    .X(_19868_));
 sky130_fd_sc_hd__buf_8 _23655_ (.A(_19868_),
    .X(_19869_));
 sky130_fd_sc_hd__buf_6 _23656_ (.A(_19869_),
    .X(_19870_));
 sky130_fd_sc_hd__mux2_1 _23657_ (.A0(_19870_),
    .A1(_19796_),
    .S(_19857_),
    .X(_03047_));
 sky130_fd_sc_hd__buf_6 _23658_ (.A(\pcpi_mul.rs1[19] ),
    .X(_19871_));
 sky130_fd_sc_hd__buf_2 _23659_ (.A(_19871_),
    .X(_19872_));
 sky130_fd_sc_hd__mux2_1 _23660_ (.A0(_19872_),
    .A1(_19797_),
    .S(_19857_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_4 _23661_ (.A(\pcpi_mul.rs1[18] ),
    .X(_19873_));
 sky130_fd_sc_hd__clkbuf_8 _23662_ (.A(_19873_),
    .X(_19874_));
 sky130_fd_sc_hd__buf_6 _23663_ (.A(_19874_),
    .X(_19875_));
 sky130_fd_sc_hd__buf_2 _23664_ (.A(_19638_),
    .X(_19876_));
 sky130_fd_sc_hd__mux2_1 _23665_ (.A0(_19875_),
    .A1(_19799_),
    .S(_19876_),
    .X(_03045_));
 sky130_fd_sc_hd__buf_6 _23666_ (.A(\pcpi_mul.rs1[17] ),
    .X(_19877_));
 sky130_fd_sc_hd__buf_6 _23667_ (.A(_19877_),
    .X(_19878_));
 sky130_fd_sc_hd__buf_6 _23668_ (.A(_19878_),
    .X(_19879_));
 sky130_fd_sc_hd__mux2_1 _23669_ (.A0(_19879_),
    .A1(_19800_),
    .S(_19876_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_4 _23670_ (.A(\pcpi_mul.rs1[16] ),
    .X(_19880_));
 sky130_fd_sc_hd__buf_6 _23671_ (.A(net497),
    .X(_19881_));
 sky130_fd_sc_hd__buf_2 _23672_ (.A(_19881_),
    .X(_19882_));
 sky130_fd_sc_hd__mux2_1 _23673_ (.A0(net454),
    .A1(_19801_),
    .S(_19876_),
    .X(_03043_));
 sky130_fd_sc_hd__buf_4 _23674_ (.A(\pcpi_mul.rs1[15] ),
    .X(_19883_));
 sky130_fd_sc_hd__buf_6 _23675_ (.A(_19883_),
    .X(_19884_));
 sky130_fd_sc_hd__clkbuf_8 _23676_ (.A(_19884_),
    .X(_19885_));
 sky130_fd_sc_hd__mux2_1 _23677_ (.A0(_19885_),
    .A1(_19802_),
    .S(_19876_),
    .X(_03042_));
 sky130_fd_sc_hd__buf_2 _23678_ (.A(\pcpi_mul.rs1[14] ),
    .X(_19886_));
 sky130_fd_sc_hd__buf_4 _23679_ (.A(_19886_),
    .X(_19887_));
 sky130_fd_sc_hd__clkbuf_4 _23680_ (.A(_19887_),
    .X(_19888_));
 sky130_fd_sc_hd__buf_1 _23681_ (.A(_19888_),
    .X(_19889_));
 sky130_fd_sc_hd__mux2_1 _23682_ (.A0(net435),
    .A1(_19803_),
    .S(_19876_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_4 _23683_ (.A(\pcpi_mul.rs1[13] ),
    .X(_19890_));
 sky130_fd_sc_hd__buf_4 _23684_ (.A(_19890_),
    .X(_19891_));
 sky130_fd_sc_hd__buf_6 _23685_ (.A(_19891_),
    .X(_19892_));
 sky130_fd_sc_hd__mux2_1 _23686_ (.A0(_19892_),
    .A1(_19804_),
    .S(_19876_),
    .X(_03040_));
 sky130_fd_sc_hd__buf_6 _23687_ (.A(\pcpi_mul.rs1[12] ),
    .X(_19893_));
 sky130_fd_sc_hd__buf_6 _23688_ (.A(_19893_),
    .X(_19894_));
 sky130_fd_sc_hd__buf_6 _23689_ (.A(_19894_),
    .X(_19895_));
 sky130_fd_sc_hd__buf_2 _23690_ (.A(_18463_),
    .X(_19896_));
 sky130_fd_sc_hd__mux2_1 _23691_ (.A0(_19895_),
    .A1(_19806_),
    .S(_19896_),
    .X(_03039_));
 sky130_fd_sc_hd__buf_4 _23692_ (.A(\pcpi_mul.rs1[11] ),
    .X(_19897_));
 sky130_fd_sc_hd__buf_6 _23693_ (.A(_19897_),
    .X(_19898_));
 sky130_fd_sc_hd__clkbuf_8 _23694_ (.A(_19898_),
    .X(_19899_));
 sky130_fd_sc_hd__mux2_1 _23695_ (.A0(_19899_),
    .A1(_19807_),
    .S(_19896_),
    .X(_03038_));
 sky130_fd_sc_hd__buf_2 _23696_ (.A(\pcpi_mul.rs1[10] ),
    .X(_19900_));
 sky130_fd_sc_hd__buf_6 _23697_ (.A(_19900_),
    .X(_19901_));
 sky130_fd_sc_hd__buf_6 _23698_ (.A(_19901_),
    .X(_19902_));
 sky130_fd_sc_hd__mux2_1 _23699_ (.A0(_19902_),
    .A1(_19808_),
    .S(_19896_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_4 _23700_ (.A(\pcpi_mul.rs1[9] ),
    .X(_19903_));
 sky130_fd_sc_hd__buf_6 _23701_ (.A(_19903_),
    .X(_19904_));
 sky130_fd_sc_hd__buf_6 _23702_ (.A(_19904_),
    .X(_19905_));
 sky130_fd_sc_hd__mux2_1 _23703_ (.A0(_19905_),
    .A1(_19809_),
    .S(_19896_),
    .X(_03036_));
 sky130_fd_sc_hd__buf_4 _23704_ (.A(\pcpi_mul.rs1[8] ),
    .X(_19906_));
 sky130_fd_sc_hd__buf_6 _23705_ (.A(_19906_),
    .X(_19907_));
 sky130_fd_sc_hd__buf_6 _23706_ (.A(_19907_),
    .X(_19908_));
 sky130_fd_sc_hd__mux2_1 _23707_ (.A0(_19908_),
    .A1(_19810_),
    .S(_19896_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_8 _23708_ (.A(\pcpi_mul.rs1[7] ),
    .X(_19909_));
 sky130_fd_sc_hd__buf_4 _23709_ (.A(_19909_),
    .X(_19910_));
 sky130_fd_sc_hd__buf_6 _23710_ (.A(_19910_),
    .X(_19911_));
 sky130_fd_sc_hd__mux2_1 _23711_ (.A0(_19911_),
    .A1(_19811_),
    .S(_19896_),
    .X(_03034_));
 sky130_fd_sc_hd__buf_4 _23712_ (.A(\pcpi_mul.rs1[6] ),
    .X(_19912_));
 sky130_fd_sc_hd__buf_4 _23713_ (.A(_19912_),
    .X(_19913_));
 sky130_fd_sc_hd__buf_6 _23714_ (.A(_19913_),
    .X(_19914_));
 sky130_fd_sc_hd__buf_2 _23715_ (.A(_18463_),
    .X(_19915_));
 sky130_fd_sc_hd__mux2_1 _23716_ (.A0(_19914_),
    .A1(_19813_),
    .S(_19915_),
    .X(_03033_));
 sky130_fd_sc_hd__buf_4 _23717_ (.A(\pcpi_mul.rs1[5] ),
    .X(_19916_));
 sky130_fd_sc_hd__buf_6 _23718_ (.A(_19916_),
    .X(_19917_));
 sky130_fd_sc_hd__buf_6 _23719_ (.A(_19917_),
    .X(_19918_));
 sky130_fd_sc_hd__mux2_1 _23720_ (.A0(_19918_),
    .A1(_19814_),
    .S(_19915_),
    .X(_03032_));
 sky130_fd_sc_hd__buf_6 _23721_ (.A(\pcpi_mul.rs1[4] ),
    .X(_19919_));
 sky130_fd_sc_hd__buf_6 _23722_ (.A(_19919_),
    .X(_19920_));
 sky130_fd_sc_hd__buf_6 _23723_ (.A(_19920_),
    .X(_19921_));
 sky130_fd_sc_hd__mux2_1 _23724_ (.A0(_19921_),
    .A1(_19815_),
    .S(_19915_),
    .X(_03031_));
 sky130_fd_sc_hd__buf_6 _23725_ (.A(\pcpi_mul.rs1[3] ),
    .X(_19922_));
 sky130_fd_sc_hd__buf_8 _23726_ (.A(_19922_),
    .X(_19923_));
 sky130_fd_sc_hd__buf_4 _23727_ (.A(_19923_),
    .X(_19924_));
 sky130_fd_sc_hd__buf_4 _23728_ (.A(_19924_),
    .X(_19925_));
 sky130_fd_sc_hd__mux2_1 _23729_ (.A0(_19925_),
    .A1(_19816_),
    .S(_19915_),
    .X(_03030_));
 sky130_fd_sc_hd__buf_6 _23730_ (.A(\pcpi_mul.rs1[2] ),
    .X(_19926_));
 sky130_fd_sc_hd__buf_6 _23731_ (.A(_19926_),
    .X(_19927_));
 sky130_fd_sc_hd__buf_4 _23732_ (.A(_19927_),
    .X(_19928_));
 sky130_fd_sc_hd__mux2_1 _23733_ (.A0(_19928_),
    .A1(_19817_),
    .S(_19915_),
    .X(_03029_));
 sky130_fd_sc_hd__buf_4 _23734_ (.A(\pcpi_mul.rs1[1] ),
    .X(_19929_));
 sky130_fd_sc_hd__clkbuf_4 _23735_ (.A(_19929_),
    .X(_19930_));
 sky130_fd_sc_hd__clkbuf_4 _23736_ (.A(_19930_),
    .X(_19931_));
 sky130_fd_sc_hd__mux2_1 _23737_ (.A0(_19931_),
    .A1(_19819_),
    .S(_19915_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_4 _23738_ (.A(\pcpi_mul.rs1[0] ),
    .X(_19932_));
 sky130_fd_sc_hd__buf_6 _23739_ (.A(_19932_),
    .X(_19933_));
 sky130_fd_sc_hd__buf_6 _23740_ (.A(_19933_),
    .X(_19934_));
 sky130_fd_sc_hd__mux2_1 _23741_ (.A0(_19934_),
    .A1(_19820_),
    .S(_18464_),
    .X(_03027_));
 sky130_fd_sc_hd__clkbuf_2 _23742_ (.A(\cpuregs_wrdata[31] ),
    .X(_19935_));
 sky130_fd_sc_hd__nand2_1 _23743_ (.A(_19415_),
    .B(_19376_),
    .Y(_19936_));
 sky130_fd_sc_hd__clkbuf_8 _23744_ (.A(_19936_),
    .X(_19937_));
 sky130_fd_sc_hd__buf_4 _23745_ (.A(_19937_),
    .X(_19938_));
 sky130_fd_sc_hd__mux2_1 _23746_ (.A0(_19935_),
    .A1(\cpuregs[5][31] ),
    .S(_19938_),
    .X(_03026_));
 sky130_fd_sc_hd__clkbuf_2 _23747_ (.A(\cpuregs_wrdata[30] ),
    .X(_19939_));
 sky130_fd_sc_hd__mux2_1 _23748_ (.A0(_19939_),
    .A1(\cpuregs[5][30] ),
    .S(_19938_),
    .X(_03025_));
 sky130_fd_sc_hd__clkbuf_2 _23749_ (.A(\cpuregs_wrdata[29] ),
    .X(_19940_));
 sky130_fd_sc_hd__mux2_1 _23750_ (.A0(_19940_),
    .A1(\cpuregs[5][29] ),
    .S(_19938_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_2 _23751_ (.A(\cpuregs_wrdata[28] ),
    .X(_19941_));
 sky130_fd_sc_hd__mux2_1 _23752_ (.A0(_19941_),
    .A1(\cpuregs[5][28] ),
    .S(_19938_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_2 _23753_ (.A(\cpuregs_wrdata[27] ),
    .X(_19942_));
 sky130_fd_sc_hd__mux2_1 _23754_ (.A0(_19942_),
    .A1(\cpuregs[5][27] ),
    .S(_19938_),
    .X(_03022_));
 sky130_fd_sc_hd__clkbuf_2 _23755_ (.A(\cpuregs_wrdata[26] ),
    .X(_19943_));
 sky130_fd_sc_hd__mux2_1 _23756_ (.A0(_19943_),
    .A1(\cpuregs[5][26] ),
    .S(_19938_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_2 _23757_ (.A(\cpuregs_wrdata[25] ),
    .X(_19944_));
 sky130_fd_sc_hd__clkbuf_4 _23758_ (.A(_19937_),
    .X(_19945_));
 sky130_fd_sc_hd__mux2_1 _23759_ (.A0(_19944_),
    .A1(\cpuregs[5][25] ),
    .S(_19945_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_2 _23760_ (.A(\cpuregs_wrdata[24] ),
    .X(_19946_));
 sky130_fd_sc_hd__mux2_1 _23761_ (.A0(_19946_),
    .A1(\cpuregs[5][24] ),
    .S(_19945_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_2 _23762_ (.A(\cpuregs_wrdata[23] ),
    .X(_19947_));
 sky130_fd_sc_hd__mux2_1 _23763_ (.A0(_19947_),
    .A1(\cpuregs[5][23] ),
    .S(_19945_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_2 _23764_ (.A(\cpuregs_wrdata[22] ),
    .X(_19948_));
 sky130_fd_sc_hd__mux2_1 _23765_ (.A0(_19948_),
    .A1(\cpuregs[5][22] ),
    .S(_19945_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_2 _23766_ (.A(\cpuregs_wrdata[21] ),
    .X(_19949_));
 sky130_fd_sc_hd__mux2_1 _23767_ (.A0(_19949_),
    .A1(\cpuregs[5][21] ),
    .S(_19945_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_2 _23768_ (.A(\cpuregs_wrdata[20] ),
    .X(_19950_));
 sky130_fd_sc_hd__mux2_1 _23769_ (.A0(_19950_),
    .A1(\cpuregs[5][20] ),
    .S(_19945_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_2 _23770_ (.A(\cpuregs_wrdata[19] ),
    .X(_19951_));
 sky130_fd_sc_hd__clkbuf_4 _23771_ (.A(_19937_),
    .X(_19952_));
 sky130_fd_sc_hd__mux2_1 _23772_ (.A0(_19951_),
    .A1(\cpuregs[5][19] ),
    .S(_19952_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_2 _23773_ (.A(\cpuregs_wrdata[18] ),
    .X(_19953_));
 sky130_fd_sc_hd__mux2_1 _23774_ (.A0(_19953_),
    .A1(\cpuregs[5][18] ),
    .S(_19952_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_2 _23775_ (.A(\cpuregs_wrdata[17] ),
    .X(_19954_));
 sky130_fd_sc_hd__mux2_1 _23776_ (.A0(_19954_),
    .A1(\cpuregs[5][17] ),
    .S(_19952_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_2 _23777_ (.A(\cpuregs_wrdata[16] ),
    .X(_19955_));
 sky130_fd_sc_hd__mux2_1 _23778_ (.A0(_19955_),
    .A1(\cpuregs[5][16] ),
    .S(_19952_),
    .X(_03011_));
 sky130_fd_sc_hd__clkbuf_2 _23779_ (.A(\cpuregs_wrdata[15] ),
    .X(_19956_));
 sky130_fd_sc_hd__mux2_1 _23780_ (.A0(_19956_),
    .A1(\cpuregs[5][15] ),
    .S(_19952_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_2 _23781_ (.A(\cpuregs_wrdata[14] ),
    .X(_19957_));
 sky130_fd_sc_hd__mux2_1 _23782_ (.A0(_19957_),
    .A1(\cpuregs[5][14] ),
    .S(_19952_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_2 _23783_ (.A(\cpuregs_wrdata[13] ),
    .X(_19958_));
 sky130_fd_sc_hd__clkbuf_4 _23784_ (.A(_19937_),
    .X(_19959_));
 sky130_fd_sc_hd__mux2_1 _23785_ (.A0(_19958_),
    .A1(\cpuregs[5][13] ),
    .S(_19959_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_2 _23786_ (.A(\cpuregs_wrdata[12] ),
    .X(_19960_));
 sky130_fd_sc_hd__mux2_1 _23787_ (.A0(_19960_),
    .A1(\cpuregs[5][12] ),
    .S(_19959_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_2 _23788_ (.A(\cpuregs_wrdata[11] ),
    .X(_19961_));
 sky130_fd_sc_hd__mux2_1 _23789_ (.A0(_19961_),
    .A1(\cpuregs[5][11] ),
    .S(_19959_),
    .X(_03006_));
 sky130_fd_sc_hd__clkbuf_2 _23790_ (.A(\cpuregs_wrdata[10] ),
    .X(_19962_));
 sky130_fd_sc_hd__mux2_1 _23791_ (.A0(_19962_),
    .A1(\cpuregs[5][10] ),
    .S(_19959_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_2 _23792_ (.A(\cpuregs_wrdata[9] ),
    .X(_19963_));
 sky130_fd_sc_hd__mux2_1 _23793_ (.A0(_19963_),
    .A1(\cpuregs[5][9] ),
    .S(_19959_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_2 _23794_ (.A(\cpuregs_wrdata[8] ),
    .X(_19964_));
 sky130_fd_sc_hd__mux2_1 _23795_ (.A0(_19964_),
    .A1(\cpuregs[5][8] ),
    .S(_19959_),
    .X(_03003_));
 sky130_fd_sc_hd__clkbuf_2 _23796_ (.A(\cpuregs_wrdata[7] ),
    .X(_19965_));
 sky130_fd_sc_hd__buf_4 _23797_ (.A(_19936_),
    .X(_19966_));
 sky130_fd_sc_hd__mux2_1 _23798_ (.A0(_19965_),
    .A1(\cpuregs[5][7] ),
    .S(_19966_),
    .X(_03002_));
 sky130_fd_sc_hd__clkbuf_2 _23799_ (.A(\cpuregs_wrdata[6] ),
    .X(_19967_));
 sky130_fd_sc_hd__mux2_1 _23800_ (.A0(_19967_),
    .A1(\cpuregs[5][6] ),
    .S(_19966_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_2 _23801_ (.A(\cpuregs_wrdata[5] ),
    .X(_19968_));
 sky130_fd_sc_hd__mux2_1 _23802_ (.A0(_19968_),
    .A1(\cpuregs[5][5] ),
    .S(_19966_),
    .X(_03000_));
 sky130_fd_sc_hd__clkbuf_2 _23803_ (.A(\cpuregs_wrdata[4] ),
    .X(_19969_));
 sky130_fd_sc_hd__mux2_1 _23804_ (.A0(_19969_),
    .A1(\cpuregs[5][4] ),
    .S(_19966_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_2 _23805_ (.A(\cpuregs_wrdata[3] ),
    .X(_19970_));
 sky130_fd_sc_hd__mux2_1 _23806_ (.A0(_19970_),
    .A1(\cpuregs[5][3] ),
    .S(_19966_),
    .X(_02998_));
 sky130_fd_sc_hd__clkbuf_2 _23807_ (.A(\cpuregs_wrdata[2] ),
    .X(_19971_));
 sky130_fd_sc_hd__mux2_1 _23808_ (.A0(_19971_),
    .A1(\cpuregs[5][2] ),
    .S(_19966_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_2 _23809_ (.A(\cpuregs_wrdata[1] ),
    .X(_19972_));
 sky130_fd_sc_hd__mux2_1 _23810_ (.A0(_19972_),
    .A1(\cpuregs[5][1] ),
    .S(_19937_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_2 _23811_ (.A(\cpuregs_wrdata[0] ),
    .X(_19973_));
 sky130_fd_sc_hd__mux2_1 _23812_ (.A0(_19973_),
    .A1(\cpuregs[5][0] ),
    .S(_19937_),
    .X(_02995_));
 sky130_fd_sc_hd__nand2_1 _23813_ (.A(_19374_),
    .B(_19538_),
    .Y(_19974_));
 sky130_fd_sc_hd__buf_8 _23814_ (.A(_19974_),
    .X(_19975_));
 sky130_fd_sc_hd__clkbuf_4 _23815_ (.A(_19975_),
    .X(_19976_));
 sky130_fd_sc_hd__mux2_1 _23816_ (.A0(_19935_),
    .A1(\cpuregs[2][31] ),
    .S(_19976_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _23817_ (.A0(_19939_),
    .A1(\cpuregs[2][30] ),
    .S(_19976_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_1 _23818_ (.A0(_19940_),
    .A1(\cpuregs[2][29] ),
    .S(_19976_),
    .X(_02992_));
 sky130_fd_sc_hd__mux2_1 _23819_ (.A0(_19941_),
    .A1(\cpuregs[2][28] ),
    .S(_19976_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _23820_ (.A0(_19942_),
    .A1(\cpuregs[2][27] ),
    .S(_19976_),
    .X(_02990_));
 sky130_fd_sc_hd__mux2_1 _23821_ (.A0(_19943_),
    .A1(\cpuregs[2][26] ),
    .S(_19976_),
    .X(_02989_));
 sky130_fd_sc_hd__buf_2 _23822_ (.A(_19975_),
    .X(_19977_));
 sky130_fd_sc_hd__mux2_1 _23823_ (.A0(_19944_),
    .A1(\cpuregs[2][25] ),
    .S(_19977_),
    .X(_02988_));
 sky130_fd_sc_hd__mux2_1 _23824_ (.A0(_19946_),
    .A1(\cpuregs[2][24] ),
    .S(_19977_),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_1 _23825_ (.A0(_19947_),
    .A1(\cpuregs[2][23] ),
    .S(_19977_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _23826_ (.A0(_19948_),
    .A1(\cpuregs[2][22] ),
    .S(_19977_),
    .X(_02985_));
 sky130_fd_sc_hd__mux2_1 _23827_ (.A0(_19949_),
    .A1(\cpuregs[2][21] ),
    .S(_19977_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2_1 _23828_ (.A0(_19950_),
    .A1(\cpuregs[2][20] ),
    .S(_19977_),
    .X(_02983_));
 sky130_fd_sc_hd__clkbuf_4 _23829_ (.A(_19975_),
    .X(_19978_));
 sky130_fd_sc_hd__mux2_1 _23830_ (.A0(_19951_),
    .A1(\cpuregs[2][19] ),
    .S(_19978_),
    .X(_02982_));
 sky130_fd_sc_hd__mux2_1 _23831_ (.A0(_19953_),
    .A1(\cpuregs[2][18] ),
    .S(_19978_),
    .X(_02981_));
 sky130_fd_sc_hd__mux2_1 _23832_ (.A0(_19954_),
    .A1(\cpuregs[2][17] ),
    .S(_19978_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _23833_ (.A0(_19955_),
    .A1(\cpuregs[2][16] ),
    .S(_19978_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _23834_ (.A0(_19956_),
    .A1(\cpuregs[2][15] ),
    .S(_19978_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_1 _23835_ (.A0(_19957_),
    .A1(\cpuregs[2][14] ),
    .S(_19978_),
    .X(_02977_));
 sky130_fd_sc_hd__buf_2 _23836_ (.A(_19975_),
    .X(_19979_));
 sky130_fd_sc_hd__mux2_1 _23837_ (.A0(_19958_),
    .A1(\cpuregs[2][13] ),
    .S(_19979_),
    .X(_02976_));
 sky130_fd_sc_hd__mux2_1 _23838_ (.A0(_19960_),
    .A1(\cpuregs[2][12] ),
    .S(_19979_),
    .X(_02975_));
 sky130_fd_sc_hd__mux2_1 _23839_ (.A0(_19961_),
    .A1(\cpuregs[2][11] ),
    .S(_19979_),
    .X(_02974_));
 sky130_fd_sc_hd__mux2_1 _23840_ (.A0(_19962_),
    .A1(\cpuregs[2][10] ),
    .S(_19979_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _23841_ (.A0(_19963_),
    .A1(\cpuregs[2][9] ),
    .S(_19979_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _23842_ (.A0(_19964_),
    .A1(\cpuregs[2][8] ),
    .S(_19979_),
    .X(_02971_));
 sky130_fd_sc_hd__buf_4 _23843_ (.A(_19974_),
    .X(_19980_));
 sky130_fd_sc_hd__mux2_1 _23844_ (.A0(_19965_),
    .A1(\cpuregs[2][7] ),
    .S(_19980_),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _23845_ (.A0(_19967_),
    .A1(\cpuregs[2][6] ),
    .S(_19980_),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _23846_ (.A0(_19968_),
    .A1(\cpuregs[2][5] ),
    .S(_19980_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _23847_ (.A0(_19969_),
    .A1(\cpuregs[2][4] ),
    .S(_19980_),
    .X(_02967_));
 sky130_fd_sc_hd__mux2_1 _23848_ (.A0(_19970_),
    .A1(\cpuregs[2][3] ),
    .S(_19980_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_1 _23849_ (.A0(_19971_),
    .A1(\cpuregs[2][2] ),
    .S(_19980_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _23850_ (.A0(_19972_),
    .A1(\cpuregs[2][1] ),
    .S(_19975_),
    .X(_02964_));
 sky130_fd_sc_hd__mux2_1 _23851_ (.A0(_19973_),
    .A1(\cpuregs[2][0] ),
    .S(_19975_),
    .X(_02963_));
 sky130_fd_sc_hd__clkbuf_4 _23852_ (.A(_18313_),
    .X(_19981_));
 sky130_fd_sc_hd__mux2_1 _23853_ (.A0(net57),
    .A1(_18672_),
    .S(_19981_),
    .X(_02962_));
 sky130_fd_sc_hd__mux2_1 _23854_ (.A0(net513),
    .A1(\mem_rdata_q[30] ),
    .S(_19981_),
    .X(_02961_));
 sky130_fd_sc_hd__mux2_1 _23855_ (.A0(net54),
    .A1(\mem_rdata_q[29] ),
    .S(_19981_),
    .X(_02960_));
 sky130_fd_sc_hd__mux2_1 _23856_ (.A0(net53),
    .A1(\mem_rdata_q[28] ),
    .S(_19981_),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_1 _23857_ (.A0(net52),
    .A1(\mem_rdata_q[27] ),
    .S(_19981_),
    .X(_02958_));
 sky130_fd_sc_hd__clkbuf_2 _23858_ (.A(_18313_),
    .X(_19982_));
 sky130_fd_sc_hd__buf_2 _23859_ (.A(_19982_),
    .X(_19983_));
 sky130_fd_sc_hd__mux2_1 _23860_ (.A0(net51),
    .A1(_19737_),
    .S(_19983_),
    .X(_02957_));
 sky130_fd_sc_hd__mux2_1 _23861_ (.A0(net50),
    .A1(\mem_rdata_q[25] ),
    .S(_19983_),
    .X(_02956_));
 sky130_fd_sc_hd__mux2_1 _23862_ (.A0(net49),
    .A1(\mem_rdata_q[24] ),
    .S(_19983_),
    .X(_02955_));
 sky130_fd_sc_hd__mux2_1 _23863_ (.A0(net48),
    .A1(\mem_rdata_q[23] ),
    .S(_19983_),
    .X(_02954_));
 sky130_fd_sc_hd__mux2_1 _23864_ (.A0(net47),
    .A1(\mem_rdata_q[22] ),
    .S(_19983_),
    .X(_02953_));
 sky130_fd_sc_hd__mux2_1 _23865_ (.A0(net46),
    .A1(\mem_rdata_q[21] ),
    .S(_19983_),
    .X(_02952_));
 sky130_fd_sc_hd__buf_2 _23866_ (.A(_19982_),
    .X(_19984_));
 sky130_fd_sc_hd__mux2_1 _23867_ (.A0(net514),
    .A1(\mem_rdata_q[20] ),
    .S(_19984_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _23868_ (.A0(net515),
    .A1(\mem_rdata_q[19] ),
    .S(_19984_),
    .X(_02950_));
 sky130_fd_sc_hd__mux2_1 _23869_ (.A0(net42),
    .A1(\mem_rdata_q[18] ),
    .S(_19984_),
    .X(_02949_));
 sky130_fd_sc_hd__mux2_1 _23870_ (.A0(net41),
    .A1(\mem_rdata_q[17] ),
    .S(_19984_),
    .X(_02948_));
 sky130_fd_sc_hd__mux2_1 _23871_ (.A0(net40),
    .A1(\mem_rdata_q[16] ),
    .S(_19984_),
    .X(_02947_));
 sky130_fd_sc_hd__mux2_1 _23872_ (.A0(net516),
    .A1(\mem_rdata_q[15] ),
    .S(_19984_),
    .X(_02946_));
 sky130_fd_sc_hd__buf_2 _23873_ (.A(_19982_),
    .X(_19985_));
 sky130_fd_sc_hd__mux2_1 _23874_ (.A0(net38),
    .A1(_18667_),
    .S(_19985_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_1 _23875_ (.A0(net37),
    .A1(\mem_rdata_q[13] ),
    .S(_19985_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _23876_ (.A0(net517),
    .A1(_18692_),
    .S(_19985_),
    .X(_02943_));
 sky130_fd_sc_hd__mux2_1 _23877_ (.A0(net35),
    .A1(\mem_rdata_q[11] ),
    .S(_19985_),
    .X(_02942_));
 sky130_fd_sc_hd__mux2_1 _23878_ (.A0(net34),
    .A1(\mem_rdata_q[10] ),
    .S(_19985_),
    .X(_02941_));
 sky130_fd_sc_hd__mux2_1 _23879_ (.A0(net64),
    .A1(\mem_rdata_q[9] ),
    .S(_19985_),
    .X(_02940_));
 sky130_fd_sc_hd__buf_2 _23880_ (.A(_18313_),
    .X(_19986_));
 sky130_fd_sc_hd__mux2_1 _23881_ (.A0(net63),
    .A1(\mem_rdata_q[8] ),
    .S(_19986_),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _23882_ (.A0(net62),
    .A1(\mem_rdata_q[7] ),
    .S(_19986_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _23883_ (.A0(net61),
    .A1(\mem_rdata_q[6] ),
    .S(_19986_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _23884_ (.A0(net512),
    .A1(\mem_rdata_q[5] ),
    .S(_19986_),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_1 _23885_ (.A0(net59),
    .A1(\mem_rdata_q[4] ),
    .S(_19986_),
    .X(_02935_));
 sky130_fd_sc_hd__mux2_1 _23886_ (.A0(net58),
    .A1(\mem_rdata_q[3] ),
    .S(_19986_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_1 _23887_ (.A0(net55),
    .A1(\mem_rdata_q[2] ),
    .S(_19982_),
    .X(_02933_));
 sky130_fd_sc_hd__mux2_1 _23888_ (.A0(net44),
    .A1(\mem_rdata_q[1] ),
    .S(_19982_),
    .X(_02932_));
 sky130_fd_sc_hd__mux2_1 _23889_ (.A0(net33),
    .A1(\mem_rdata_q[0] ),
    .S(_19982_),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_1 _23890_ (.A(_19374_),
    .B(_19464_),
    .Y(_19987_));
 sky130_fd_sc_hd__buf_6 _23891_ (.A(_19987_),
    .X(_19988_));
 sky130_fd_sc_hd__clkbuf_4 _23892_ (.A(_19988_),
    .X(_19989_));
 sky130_fd_sc_hd__mux2_1 _23893_ (.A0(_19935_),
    .A1(\cpuregs[18][31] ),
    .S(_19989_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _23894_ (.A0(_19939_),
    .A1(\cpuregs[18][30] ),
    .S(_19989_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_1 _23895_ (.A0(_19940_),
    .A1(\cpuregs[18][29] ),
    .S(_19989_),
    .X(_02928_));
 sky130_fd_sc_hd__mux2_1 _23896_ (.A0(_19941_),
    .A1(\cpuregs[18][28] ),
    .S(_19989_),
    .X(_02927_));
 sky130_fd_sc_hd__mux2_1 _23897_ (.A0(_19942_),
    .A1(\cpuregs[18][27] ),
    .S(_19989_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _23898_ (.A0(_19943_),
    .A1(\cpuregs[18][26] ),
    .S(_19989_),
    .X(_02925_));
 sky130_fd_sc_hd__clkbuf_4 _23899_ (.A(_19988_),
    .X(_19990_));
 sky130_fd_sc_hd__mux2_1 _23900_ (.A0(_19944_),
    .A1(\cpuregs[18][25] ),
    .S(_19990_),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_1 _23901_ (.A0(_19946_),
    .A1(\cpuregs[18][24] ),
    .S(_19990_),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _23902_ (.A0(_19947_),
    .A1(\cpuregs[18][23] ),
    .S(_19990_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _23903_ (.A0(_19948_),
    .A1(\cpuregs[18][22] ),
    .S(_19990_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _23904_ (.A0(_19949_),
    .A1(\cpuregs[18][21] ),
    .S(_19990_),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_1 _23905_ (.A0(_19950_),
    .A1(\cpuregs[18][20] ),
    .S(_19990_),
    .X(_02919_));
 sky130_fd_sc_hd__clkbuf_4 _23906_ (.A(_19988_),
    .X(_19991_));
 sky130_fd_sc_hd__mux2_1 _23907_ (.A0(_19951_),
    .A1(\cpuregs[18][19] ),
    .S(_19991_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _23908_ (.A0(_19953_),
    .A1(\cpuregs[18][18] ),
    .S(_19991_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _23909_ (.A0(_19954_),
    .A1(\cpuregs[18][17] ),
    .S(_19991_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _23910_ (.A0(_19955_),
    .A1(\cpuregs[18][16] ),
    .S(_19991_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _23911_ (.A0(_19956_),
    .A1(\cpuregs[18][15] ),
    .S(_19991_),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _23912_ (.A0(_19957_),
    .A1(\cpuregs[18][14] ),
    .S(_19991_),
    .X(_02913_));
 sky130_fd_sc_hd__buf_2 _23913_ (.A(_19988_),
    .X(_19992_));
 sky130_fd_sc_hd__mux2_1 _23914_ (.A0(_19958_),
    .A1(\cpuregs[18][13] ),
    .S(_19992_),
    .X(_02912_));
 sky130_fd_sc_hd__mux2_1 _23915_ (.A0(_19960_),
    .A1(\cpuregs[18][12] ),
    .S(_19992_),
    .X(_02911_));
 sky130_fd_sc_hd__mux2_1 _23916_ (.A0(_19961_),
    .A1(\cpuregs[18][11] ),
    .S(_19992_),
    .X(_02910_));
 sky130_fd_sc_hd__mux2_1 _23917_ (.A0(_19962_),
    .A1(\cpuregs[18][10] ),
    .S(_19992_),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_1 _23918_ (.A0(_19963_),
    .A1(\cpuregs[18][9] ),
    .S(_19992_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _23919_ (.A0(_19964_),
    .A1(\cpuregs[18][8] ),
    .S(_19992_),
    .X(_02907_));
 sky130_fd_sc_hd__clkbuf_4 _23920_ (.A(_19987_),
    .X(_19993_));
 sky130_fd_sc_hd__mux2_1 _23921_ (.A0(_19965_),
    .A1(\cpuregs[18][7] ),
    .S(_19993_),
    .X(_02906_));
 sky130_fd_sc_hd__mux2_1 _23922_ (.A0(_19967_),
    .A1(\cpuregs[18][6] ),
    .S(_19993_),
    .X(_02905_));
 sky130_fd_sc_hd__mux2_1 _23923_ (.A0(_19968_),
    .A1(\cpuregs[18][5] ),
    .S(_19993_),
    .X(_02904_));
 sky130_fd_sc_hd__mux2_1 _23924_ (.A0(_19969_),
    .A1(\cpuregs[18][4] ),
    .S(_19993_),
    .X(_02903_));
 sky130_fd_sc_hd__mux2_1 _23925_ (.A0(_19970_),
    .A1(\cpuregs[18][3] ),
    .S(_19993_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_1 _23926_ (.A0(_19971_),
    .A1(\cpuregs[18][2] ),
    .S(_19993_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _23927_ (.A0(_19972_),
    .A1(\cpuregs[18][1] ),
    .S(_19988_),
    .X(_02900_));
 sky130_fd_sc_hd__mux2_1 _23928_ (.A0(_19973_),
    .A1(\cpuregs[18][0] ),
    .S(_19988_),
    .X(_02899_));
 sky130_fd_sc_hd__nand2_1 _23929_ (.A(_19374_),
    .B(_19417_),
    .Y(_19994_));
 sky130_fd_sc_hd__clkbuf_8 _23930_ (.A(_19994_),
    .X(_19995_));
 sky130_fd_sc_hd__buf_4 _23931_ (.A(_19995_),
    .X(_19996_));
 sky130_fd_sc_hd__mux2_1 _23932_ (.A0(_19935_),
    .A1(\cpuregs[10][31] ),
    .S(_19996_),
    .X(_02898_));
 sky130_fd_sc_hd__mux2_1 _23933_ (.A0(_19939_),
    .A1(\cpuregs[10][30] ),
    .S(_19996_),
    .X(_02897_));
 sky130_fd_sc_hd__mux2_1 _23934_ (.A0(_19940_),
    .A1(\cpuregs[10][29] ),
    .S(_19996_),
    .X(_02896_));
 sky130_fd_sc_hd__mux2_1 _23935_ (.A0(_19941_),
    .A1(\cpuregs[10][28] ),
    .S(_19996_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _23936_ (.A0(_19942_),
    .A1(\cpuregs[10][27] ),
    .S(_19996_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _23937_ (.A0(_19943_),
    .A1(\cpuregs[10][26] ),
    .S(_19996_),
    .X(_02893_));
 sky130_fd_sc_hd__buf_2 _23938_ (.A(_19995_),
    .X(_19997_));
 sky130_fd_sc_hd__mux2_1 _23939_ (.A0(_19944_),
    .A1(\cpuregs[10][25] ),
    .S(_19997_),
    .X(_02892_));
 sky130_fd_sc_hd__mux2_1 _23940_ (.A0(_19946_),
    .A1(\cpuregs[10][24] ),
    .S(_19997_),
    .X(_02891_));
 sky130_fd_sc_hd__mux2_1 _23941_ (.A0(_19947_),
    .A1(\cpuregs[10][23] ),
    .S(_19997_),
    .X(_02890_));
 sky130_fd_sc_hd__mux2_1 _23942_ (.A0(_19948_),
    .A1(\cpuregs[10][22] ),
    .S(_19997_),
    .X(_02889_));
 sky130_fd_sc_hd__mux2_1 _23943_ (.A0(_19949_),
    .A1(\cpuregs[10][21] ),
    .S(_19997_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _23944_ (.A0(_19950_),
    .A1(\cpuregs[10][20] ),
    .S(_19997_),
    .X(_02887_));
 sky130_fd_sc_hd__clkbuf_4 _23945_ (.A(_19995_),
    .X(_19998_));
 sky130_fd_sc_hd__mux2_1 _23946_ (.A0(_19951_),
    .A1(\cpuregs[10][19] ),
    .S(_19998_),
    .X(_02886_));
 sky130_fd_sc_hd__mux2_1 _23947_ (.A0(_19953_),
    .A1(\cpuregs[10][18] ),
    .S(_19998_),
    .X(_02885_));
 sky130_fd_sc_hd__mux2_1 _23948_ (.A0(_19954_),
    .A1(\cpuregs[10][17] ),
    .S(_19998_),
    .X(_02884_));
 sky130_fd_sc_hd__mux2_1 _23949_ (.A0(_19955_),
    .A1(\cpuregs[10][16] ),
    .S(_19998_),
    .X(_02883_));
 sky130_fd_sc_hd__mux2_1 _23950_ (.A0(_19956_),
    .A1(\cpuregs[10][15] ),
    .S(_19998_),
    .X(_02882_));
 sky130_fd_sc_hd__mux2_1 _23951_ (.A0(_19957_),
    .A1(\cpuregs[10][14] ),
    .S(_19998_),
    .X(_02881_));
 sky130_fd_sc_hd__clkbuf_4 _23952_ (.A(_19995_),
    .X(_19999_));
 sky130_fd_sc_hd__mux2_1 _23953_ (.A0(_19958_),
    .A1(\cpuregs[10][13] ),
    .S(_19999_),
    .X(_02880_));
 sky130_fd_sc_hd__mux2_1 _23954_ (.A0(_19960_),
    .A1(\cpuregs[10][12] ),
    .S(_19999_),
    .X(_02879_));
 sky130_fd_sc_hd__mux2_1 _23955_ (.A0(_19961_),
    .A1(\cpuregs[10][11] ),
    .S(_19999_),
    .X(_02878_));
 sky130_fd_sc_hd__mux2_1 _23956_ (.A0(_19962_),
    .A1(\cpuregs[10][10] ),
    .S(_19999_),
    .X(_02877_));
 sky130_fd_sc_hd__mux2_1 _23957_ (.A0(_19963_),
    .A1(\cpuregs[10][9] ),
    .S(_19999_),
    .X(_02876_));
 sky130_fd_sc_hd__mux2_1 _23958_ (.A0(_19964_),
    .A1(\cpuregs[10][8] ),
    .S(_19999_),
    .X(_02875_));
 sky130_fd_sc_hd__buf_4 _23959_ (.A(_19994_),
    .X(_20000_));
 sky130_fd_sc_hd__mux2_1 _23960_ (.A0(_19965_),
    .A1(\cpuregs[10][7] ),
    .S(_20000_),
    .X(_02874_));
 sky130_fd_sc_hd__mux2_1 _23961_ (.A0(_19967_),
    .A1(\cpuregs[10][6] ),
    .S(_20000_),
    .X(_02873_));
 sky130_fd_sc_hd__mux2_1 _23962_ (.A0(_19968_),
    .A1(\cpuregs[10][5] ),
    .S(_20000_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _23963_ (.A0(_19969_),
    .A1(\cpuregs[10][4] ),
    .S(_20000_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _23964_ (.A0(_19970_),
    .A1(\cpuregs[10][3] ),
    .S(_20000_),
    .X(_02870_));
 sky130_fd_sc_hd__mux2_1 _23965_ (.A0(_19971_),
    .A1(\cpuregs[10][2] ),
    .S(_20000_),
    .X(_02869_));
 sky130_fd_sc_hd__mux2_1 _23966_ (.A0(_19972_),
    .A1(\cpuregs[10][1] ),
    .S(_19995_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _23967_ (.A0(_19973_),
    .A1(\cpuregs[10][0] ),
    .S(_19995_),
    .X(_02867_));
 sky130_fd_sc_hd__clkbuf_1 _23968_ (.A(\cpuregs[0][31] ),
    .X(_02866_));
 sky130_fd_sc_hd__clkbuf_1 _23969_ (.A(\cpuregs[0][30] ),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _23970_ (.A(\cpuregs[0][29] ),
    .X(_02864_));
 sky130_fd_sc_hd__clkbuf_1 _23971_ (.A(\cpuregs[0][28] ),
    .X(_02863_));
 sky130_fd_sc_hd__clkbuf_1 _23972_ (.A(\cpuregs[0][27] ),
    .X(_02862_));
 sky130_fd_sc_hd__clkbuf_1 _23973_ (.A(\cpuregs[0][26] ),
    .X(_02861_));
 sky130_fd_sc_hd__clkbuf_1 _23974_ (.A(\cpuregs[0][25] ),
    .X(_02860_));
 sky130_fd_sc_hd__clkbuf_1 _23975_ (.A(\cpuregs[0][24] ),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _23976_ (.A(\cpuregs[0][23] ),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_1 _23977_ (.A(\cpuregs[0][22] ),
    .X(_02857_));
 sky130_fd_sc_hd__clkbuf_1 _23978_ (.A(\cpuregs[0][21] ),
    .X(_02856_));
 sky130_fd_sc_hd__clkbuf_1 _23979_ (.A(\cpuregs[0][20] ),
    .X(_02855_));
 sky130_fd_sc_hd__clkbuf_1 _23980_ (.A(\cpuregs[0][19] ),
    .X(_02854_));
 sky130_fd_sc_hd__clkbuf_1 _23981_ (.A(\cpuregs[0][18] ),
    .X(_02853_));
 sky130_fd_sc_hd__clkbuf_1 _23982_ (.A(\cpuregs[0][17] ),
    .X(_02852_));
 sky130_fd_sc_hd__clkbuf_1 _23983_ (.A(\cpuregs[0][16] ),
    .X(_02851_));
 sky130_fd_sc_hd__clkbuf_1 _23984_ (.A(\cpuregs[0][15] ),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _23985_ (.A(\cpuregs[0][14] ),
    .X(_02849_));
 sky130_fd_sc_hd__clkbuf_1 _23986_ (.A(\cpuregs[0][13] ),
    .X(_02848_));
 sky130_fd_sc_hd__clkbuf_1 _23987_ (.A(\cpuregs[0][12] ),
    .X(_02847_));
 sky130_fd_sc_hd__clkbuf_1 _23988_ (.A(\cpuregs[0][11] ),
    .X(_02846_));
 sky130_fd_sc_hd__clkbuf_1 _23989_ (.A(\cpuregs[0][10] ),
    .X(_02845_));
 sky130_fd_sc_hd__clkbuf_1 _23990_ (.A(\cpuregs[0][9] ),
    .X(_02844_));
 sky130_fd_sc_hd__clkbuf_1 _23991_ (.A(\cpuregs[0][8] ),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _23992_ (.A(\cpuregs[0][7] ),
    .X(_02842_));
 sky130_fd_sc_hd__clkbuf_1 _23993_ (.A(\cpuregs[0][6] ),
    .X(_02841_));
 sky130_fd_sc_hd__clkbuf_1 _23994_ (.A(\cpuregs[0][5] ),
    .X(_02840_));
 sky130_fd_sc_hd__clkbuf_1 _23995_ (.A(\cpuregs[0][4] ),
    .X(_02839_));
 sky130_fd_sc_hd__clkbuf_1 _23996_ (.A(\cpuregs[0][3] ),
    .X(_02838_));
 sky130_fd_sc_hd__clkbuf_1 _23997_ (.A(\cpuregs[0][2] ),
    .X(_02837_));
 sky130_fd_sc_hd__clkbuf_1 _23998_ (.A(\cpuregs[0][1] ),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _23999_ (.A(\cpuregs[0][0] ),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_1 _24000_ (.A(_19374_),
    .B(_19491_),
    .Y(_20001_));
 sky130_fd_sc_hd__buf_8 _24001_ (.A(_20001_),
    .X(_20002_));
 sky130_fd_sc_hd__clkbuf_4 _24002_ (.A(_20002_),
    .X(_20003_));
 sky130_fd_sc_hd__mux2_1 _24003_ (.A0(_19935_),
    .A1(\cpuregs[14][31] ),
    .S(_20003_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _24004_ (.A0(_19939_),
    .A1(\cpuregs[14][30] ),
    .S(_20003_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _24005_ (.A0(_19940_),
    .A1(\cpuregs[14][29] ),
    .S(_20003_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _24006_ (.A0(_19941_),
    .A1(\cpuregs[14][28] ),
    .S(_20003_),
    .X(_02831_));
 sky130_fd_sc_hd__mux2_1 _24007_ (.A0(_19942_),
    .A1(\cpuregs[14][27] ),
    .S(_20003_),
    .X(_02830_));
 sky130_fd_sc_hd__mux2_1 _24008_ (.A0(_19943_),
    .A1(\cpuregs[14][26] ),
    .S(_20003_),
    .X(_02829_));
 sky130_fd_sc_hd__buf_2 _24009_ (.A(_20002_),
    .X(_20004_));
 sky130_fd_sc_hd__mux2_1 _24010_ (.A0(_19944_),
    .A1(\cpuregs[14][25] ),
    .S(_20004_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _24011_ (.A0(_19946_),
    .A1(\cpuregs[14][24] ),
    .S(_20004_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _24012_ (.A0(_19947_),
    .A1(\cpuregs[14][23] ),
    .S(_20004_),
    .X(_02826_));
 sky130_fd_sc_hd__mux2_1 _24013_ (.A0(_19948_),
    .A1(\cpuregs[14][22] ),
    .S(_20004_),
    .X(_02825_));
 sky130_fd_sc_hd__mux2_1 _24014_ (.A0(_19949_),
    .A1(\cpuregs[14][21] ),
    .S(_20004_),
    .X(_02824_));
 sky130_fd_sc_hd__mux2_1 _24015_ (.A0(_19950_),
    .A1(\cpuregs[14][20] ),
    .S(_20004_),
    .X(_02823_));
 sky130_fd_sc_hd__clkbuf_4 _24016_ (.A(_20002_),
    .X(_20005_));
 sky130_fd_sc_hd__mux2_1 _24017_ (.A0(_19951_),
    .A1(\cpuregs[14][19] ),
    .S(_20005_),
    .X(_02822_));
 sky130_fd_sc_hd__mux2_1 _24018_ (.A0(_19953_),
    .A1(\cpuregs[14][18] ),
    .S(_20005_),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_1 _24019_ (.A0(_19954_),
    .A1(\cpuregs[14][17] ),
    .S(_20005_),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_1 _24020_ (.A0(_19955_),
    .A1(\cpuregs[14][16] ),
    .S(_20005_),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_1 _24021_ (.A0(_19956_),
    .A1(\cpuregs[14][15] ),
    .S(_20005_),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _24022_ (.A0(_19957_),
    .A1(\cpuregs[14][14] ),
    .S(_20005_),
    .X(_02817_));
 sky130_fd_sc_hd__buf_2 _24023_ (.A(_20002_),
    .X(_20006_));
 sky130_fd_sc_hd__mux2_1 _24024_ (.A0(_19958_),
    .A1(\cpuregs[14][13] ),
    .S(_20006_),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _24025_ (.A0(_19960_),
    .A1(\cpuregs[14][12] ),
    .S(_20006_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _24026_ (.A0(_19961_),
    .A1(\cpuregs[14][11] ),
    .S(_20006_),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _24027_ (.A0(_19962_),
    .A1(\cpuregs[14][10] ),
    .S(_20006_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _24028_ (.A0(_19963_),
    .A1(\cpuregs[14][9] ),
    .S(_20006_),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _24029_ (.A0(_19964_),
    .A1(\cpuregs[14][8] ),
    .S(_20006_),
    .X(_02811_));
 sky130_fd_sc_hd__clkbuf_4 _24030_ (.A(_20001_),
    .X(_20007_));
 sky130_fd_sc_hd__mux2_1 _24031_ (.A0(_19965_),
    .A1(\cpuregs[14][7] ),
    .S(_20007_),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _24032_ (.A0(_19967_),
    .A1(\cpuregs[14][6] ),
    .S(_20007_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _24033_ (.A0(_19968_),
    .A1(\cpuregs[14][5] ),
    .S(_20007_),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _24034_ (.A0(_19969_),
    .A1(\cpuregs[14][4] ),
    .S(_20007_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _24035_ (.A0(_19970_),
    .A1(\cpuregs[14][3] ),
    .S(_20007_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _24036_ (.A0(_19971_),
    .A1(\cpuregs[14][2] ),
    .S(_20007_),
    .X(_02805_));
 sky130_fd_sc_hd__mux2_1 _24037_ (.A0(_19972_),
    .A1(\cpuregs[14][1] ),
    .S(_20002_),
    .X(_02804_));
 sky130_fd_sc_hd__mux2_1 _24038_ (.A0(_19973_),
    .A1(\cpuregs[14][0] ),
    .S(_20002_),
    .X(_02803_));
 sky130_fd_sc_hd__or3_4 _24039_ (.A(_19366_),
    .B(_19416_),
    .C(_19372_),
    .X(_20008_));
 sky130_fd_sc_hd__clkbuf_8 _24040_ (.A(_20008_),
    .X(_20009_));
 sky130_fd_sc_hd__clkbuf_4 _24041_ (.A(_20009_),
    .X(_20010_));
 sky130_fd_sc_hd__mux2_1 _24042_ (.A0(_19935_),
    .A1(\cpuregs[8][31] ),
    .S(_20010_),
    .X(_02802_));
 sky130_fd_sc_hd__mux2_1 _24043_ (.A0(_19939_),
    .A1(\cpuregs[8][30] ),
    .S(_20010_),
    .X(_02801_));
 sky130_fd_sc_hd__mux2_1 _24044_ (.A0(_19940_),
    .A1(\cpuregs[8][29] ),
    .S(_20010_),
    .X(_02800_));
 sky130_fd_sc_hd__mux2_1 _24045_ (.A0(_19941_),
    .A1(\cpuregs[8][28] ),
    .S(_20010_),
    .X(_02799_));
 sky130_fd_sc_hd__mux2_1 _24046_ (.A0(_19942_),
    .A1(\cpuregs[8][27] ),
    .S(_20010_),
    .X(_02798_));
 sky130_fd_sc_hd__mux2_1 _24047_ (.A0(_19943_),
    .A1(\cpuregs[8][26] ),
    .S(_20010_),
    .X(_02797_));
 sky130_fd_sc_hd__buf_2 _24048_ (.A(_20009_),
    .X(_20011_));
 sky130_fd_sc_hd__mux2_1 _24049_ (.A0(_19944_),
    .A1(\cpuregs[8][25] ),
    .S(_20011_),
    .X(_02796_));
 sky130_fd_sc_hd__mux2_1 _24050_ (.A0(_19946_),
    .A1(\cpuregs[8][24] ),
    .S(_20011_),
    .X(_02795_));
 sky130_fd_sc_hd__mux2_1 _24051_ (.A0(_19947_),
    .A1(\cpuregs[8][23] ),
    .S(_20011_),
    .X(_02794_));
 sky130_fd_sc_hd__mux2_1 _24052_ (.A0(_19948_),
    .A1(\cpuregs[8][22] ),
    .S(_20011_),
    .X(_02793_));
 sky130_fd_sc_hd__mux2_1 _24053_ (.A0(_19949_),
    .A1(\cpuregs[8][21] ),
    .S(_20011_),
    .X(_02792_));
 sky130_fd_sc_hd__mux2_1 _24054_ (.A0(_19950_),
    .A1(\cpuregs[8][20] ),
    .S(_20011_),
    .X(_02791_));
 sky130_fd_sc_hd__clkbuf_4 _24055_ (.A(_20009_),
    .X(_20012_));
 sky130_fd_sc_hd__mux2_1 _24056_ (.A0(_19951_),
    .A1(\cpuregs[8][19] ),
    .S(_20012_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _24057_ (.A0(_19953_),
    .A1(\cpuregs[8][18] ),
    .S(_20012_),
    .X(_02789_));
 sky130_fd_sc_hd__mux2_1 _24058_ (.A0(_19954_),
    .A1(\cpuregs[8][17] ),
    .S(_20012_),
    .X(_02788_));
 sky130_fd_sc_hd__mux2_1 _24059_ (.A0(_19955_),
    .A1(\cpuregs[8][16] ),
    .S(_20012_),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _24060_ (.A0(_19956_),
    .A1(\cpuregs[8][15] ),
    .S(_20012_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _24061_ (.A0(_19957_),
    .A1(\cpuregs[8][14] ),
    .S(_20012_),
    .X(_02785_));
 sky130_fd_sc_hd__buf_2 _24062_ (.A(_20009_),
    .X(_20013_));
 sky130_fd_sc_hd__mux2_1 _24063_ (.A0(_19958_),
    .A1(\cpuregs[8][13] ),
    .S(_20013_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _24064_ (.A0(_19960_),
    .A1(\cpuregs[8][12] ),
    .S(_20013_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _24065_ (.A0(_19961_),
    .A1(\cpuregs[8][11] ),
    .S(_20013_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _24066_ (.A0(_19962_),
    .A1(\cpuregs[8][10] ),
    .S(_20013_),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _24067_ (.A0(_19963_),
    .A1(\cpuregs[8][9] ),
    .S(_20013_),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_1 _24068_ (.A0(_19964_),
    .A1(\cpuregs[8][8] ),
    .S(_20013_),
    .X(_02779_));
 sky130_fd_sc_hd__clkbuf_4 _24069_ (.A(_20008_),
    .X(_20014_));
 sky130_fd_sc_hd__mux2_1 _24070_ (.A0(_19965_),
    .A1(\cpuregs[8][7] ),
    .S(_20014_),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _24071_ (.A0(_19967_),
    .A1(\cpuregs[8][6] ),
    .S(_20014_),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _24072_ (.A0(_19968_),
    .A1(\cpuregs[8][5] ),
    .S(_20014_),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_1 _24073_ (.A0(_19969_),
    .A1(\cpuregs[8][4] ),
    .S(_20014_),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _24074_ (.A0(_19970_),
    .A1(\cpuregs[8][3] ),
    .S(_20014_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _24075_ (.A0(_19971_),
    .A1(\cpuregs[8][2] ),
    .S(_20014_),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _24076_ (.A0(_19972_),
    .A1(\cpuregs[8][1] ),
    .S(_20009_),
    .X(_02772_));
 sky130_fd_sc_hd__mux2_1 _24077_ (.A0(_19973_),
    .A1(\cpuregs[8][0] ),
    .S(_20009_),
    .X(_02771_));
 sky130_fd_sc_hd__nor2_8 _24078_ (.A(latched_branch),
    .B(_18525_),
    .Y(_00292_));
 sky130_fd_sc_hd__nor2_1 _24079_ (.A(_18486_),
    .B(_18344_),
    .Y(_20015_));
 sky130_fd_sc_hd__o311a_1 _24080_ (.A1(_18788_),
    .A2(_00292_),
    .A3(_20015_),
    .B1(_18333_),
    .C1(\reg_next_pc[0] ),
    .X(_02770_));
 sky130_fd_sc_hd__and2_1 _24081_ (.A(_19174_),
    .B(_00008_),
    .X(_02769_));
 sky130_fd_sc_hd__clkbuf_2 _24082_ (.A(_19173_),
    .X(_20016_));
 sky130_fd_sc_hd__and2_1 _24083_ (.A(_20016_),
    .B(_20930_),
    .X(_02768_));
 sky130_fd_sc_hd__and2_1 _24084_ (.A(_20016_),
    .B(_00031_),
    .X(_02767_));
 sky130_fd_sc_hd__and2_1 _24085_ (.A(_20016_),
    .B(_00032_),
    .X(_02766_));
 sky130_fd_sc_hd__and2_1 _24086_ (.A(_20016_),
    .B(_00033_),
    .X(_02765_));
 sky130_fd_sc_hd__and2_1 _24087_ (.A(_20016_),
    .B(_00034_),
    .X(_02764_));
 sky130_fd_sc_hd__and2_1 _24088_ (.A(_20016_),
    .B(_00035_),
    .X(_02763_));
 sky130_fd_sc_hd__clkbuf_2 _24089_ (.A(_19173_),
    .X(_20017_));
 sky130_fd_sc_hd__and2_1 _24090_ (.A(_20017_),
    .B(_00036_),
    .X(_02762_));
 sky130_fd_sc_hd__and2_1 _24091_ (.A(_20017_),
    .B(_00037_),
    .X(_02761_));
 sky130_fd_sc_hd__and2_1 _24092_ (.A(_20017_),
    .B(_00009_),
    .X(_02760_));
 sky130_fd_sc_hd__and2_1 _24093_ (.A(_20017_),
    .B(_00010_),
    .X(_02759_));
 sky130_fd_sc_hd__and2_1 _24094_ (.A(_20017_),
    .B(_00011_),
    .X(_02758_));
 sky130_fd_sc_hd__and2_1 _24095_ (.A(_20017_),
    .B(_00012_),
    .X(_02757_));
 sky130_fd_sc_hd__clkbuf_2 _24096_ (.A(_19173_),
    .X(_20018_));
 sky130_fd_sc_hd__and2_1 _24097_ (.A(_20018_),
    .B(_00013_),
    .X(_02756_));
 sky130_fd_sc_hd__and2_1 _24098_ (.A(_20018_),
    .B(_00014_),
    .X(_02755_));
 sky130_fd_sc_hd__and2_1 _24099_ (.A(_20018_),
    .B(_00015_),
    .X(_02754_));
 sky130_fd_sc_hd__and2_1 _24100_ (.A(_20018_),
    .B(_00016_),
    .X(_02753_));
 sky130_fd_sc_hd__and2_1 _24101_ (.A(_20018_),
    .B(_00017_),
    .X(_02752_));
 sky130_fd_sc_hd__and2_1 _24102_ (.A(_20018_),
    .B(_00018_),
    .X(_02751_));
 sky130_fd_sc_hd__clkbuf_2 _24103_ (.A(_19173_),
    .X(_20019_));
 sky130_fd_sc_hd__and2_1 _24104_ (.A(_20019_),
    .B(_00019_),
    .X(_02750_));
 sky130_fd_sc_hd__and2_1 _24105_ (.A(_20019_),
    .B(_00020_),
    .X(_02749_));
 sky130_fd_sc_hd__and2_1 _24106_ (.A(_20019_),
    .B(_00021_),
    .X(_02748_));
 sky130_fd_sc_hd__and2_1 _24107_ (.A(_20019_),
    .B(_00022_),
    .X(_02747_));
 sky130_fd_sc_hd__and2_1 _24108_ (.A(_20019_),
    .B(_00023_),
    .X(_02746_));
 sky130_fd_sc_hd__and2_1 _24109_ (.A(_20019_),
    .B(_00024_),
    .X(_02745_));
 sky130_fd_sc_hd__clkbuf_2 _24110_ (.A(_19173_),
    .X(_20020_));
 sky130_fd_sc_hd__and2_1 _24111_ (.A(_20020_),
    .B(_00025_),
    .X(_02744_));
 sky130_fd_sc_hd__and2_1 _24112_ (.A(_20020_),
    .B(_00026_),
    .X(_02743_));
 sky130_fd_sc_hd__and2_1 _24113_ (.A(_20020_),
    .B(_00027_),
    .X(_02742_));
 sky130_fd_sc_hd__and2_1 _24114_ (.A(_20020_),
    .B(_00028_),
    .X(_02741_));
 sky130_fd_sc_hd__and2_1 _24115_ (.A(_20020_),
    .B(_00029_),
    .X(_02740_));
 sky130_fd_sc_hd__and2_1 _24116_ (.A(_20020_),
    .B(_00030_),
    .X(_02739_));
 sky130_fd_sc_hd__or2_1 _24117_ (.A(_19764_),
    .B(_19722_),
    .X(_20021_));
 sky130_fd_sc_hd__buf_2 _24118_ (.A(instr_jal),
    .X(_20022_));
 sky130_fd_sc_hd__clkbuf_2 _24119_ (.A(_20022_),
    .X(_20023_));
 sky130_fd_sc_hd__nand2_1 _24120_ (.A(\decoded_imm_uj[1] ),
    .B(_20023_),
    .Y(_20024_));
 sky130_fd_sc_hd__nor2_2 _24121_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(is_sb_sh_sw),
    .Y(_20025_));
 sky130_vsdinv _24122_ (.A(_20025_),
    .Y(_20026_));
 sky130_fd_sc_hd__nand2_1 _24123_ (.A(_20026_),
    .B(\mem_rdata_q[8] ),
    .Y(_20027_));
 sky130_fd_sc_hd__a31o_1 _24124_ (.A1(_20021_),
    .A2(_20024_),
    .A3(_20027_),
    .B1(_18648_),
    .X(_20028_));
 sky130_fd_sc_hd__a21bo_1 _24125_ (.A1(\decoded_imm[1] ),
    .A2(_19708_),
    .B1_N(_20028_),
    .X(_02738_));
 sky130_vsdinv _24126_ (.A(\decoded_imm[2] ),
    .Y(_20029_));
 sky130_fd_sc_hd__or2b_1 _24127_ (.A(_19723_),
    .B_N(\mem_rdata_q[22] ),
    .X(_20030_));
 sky130_fd_sc_hd__clkbuf_2 _24128_ (.A(_20022_),
    .X(_20031_));
 sky130_fd_sc_hd__nand2_1 _24129_ (.A(\decoded_imm_uj[2] ),
    .B(_20031_),
    .Y(_20032_));
 sky130_fd_sc_hd__nand2_1 _24130_ (.A(_20026_),
    .B(\mem_rdata_q[9] ),
    .Y(_20033_));
 sky130_fd_sc_hd__buf_2 _24131_ (.A(_18647_),
    .X(_20034_));
 sky130_fd_sc_hd__a31o_1 _24132_ (.A1(_20030_),
    .A2(_20032_),
    .A3(_20033_),
    .B1(_20034_),
    .X(_20035_));
 sky130_fd_sc_hd__o21ai_1 _24133_ (.A1(_20029_),
    .A2(_19777_),
    .B1(_20035_),
    .Y(_02737_));
 sky130_vsdinv _24134_ (.A(\decoded_imm[3] ),
    .Y(_20036_));
 sky130_fd_sc_hd__or2b_1 _24135_ (.A(_19723_),
    .B_N(\mem_rdata_q[23] ),
    .X(_20037_));
 sky130_fd_sc_hd__nand2_1 _24136_ (.A(\decoded_imm_uj[3] ),
    .B(_20031_),
    .Y(_20038_));
 sky130_fd_sc_hd__nand2_1 _24137_ (.A(_20026_),
    .B(\mem_rdata_q[10] ),
    .Y(_20039_));
 sky130_fd_sc_hd__a31o_1 _24138_ (.A1(_20037_),
    .A2(_20038_),
    .A3(_20039_),
    .B1(_20034_),
    .X(_20040_));
 sky130_fd_sc_hd__o21ai_1 _24139_ (.A1(_20036_),
    .A2(_19777_),
    .B1(_20040_),
    .Y(_02736_));
 sky130_vsdinv _24140_ (.A(\decoded_imm[4] ),
    .Y(_20041_));
 sky130_fd_sc_hd__or2b_1 _24141_ (.A(_19723_),
    .B_N(\mem_rdata_q[24] ),
    .X(_20042_));
 sky130_fd_sc_hd__nand2_1 _24142_ (.A(\decoded_imm_uj[4] ),
    .B(_20031_),
    .Y(_20043_));
 sky130_fd_sc_hd__nand2_1 _24143_ (.A(_20026_),
    .B(\mem_rdata_q[11] ),
    .Y(_20044_));
 sky130_fd_sc_hd__a31o_1 _24144_ (.A1(_20042_),
    .A2(_20043_),
    .A3(_20044_),
    .B1(_18648_),
    .X(_20045_));
 sky130_fd_sc_hd__o21ai_1 _24145_ (.A1(_20041_),
    .A2(_19777_),
    .B1(_20045_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand2_1 _24146_ (.A(_19722_),
    .B(_20025_),
    .Y(_20046_));
 sky130_fd_sc_hd__clkbuf_2 _24147_ (.A(_20046_),
    .X(_20047_));
 sky130_fd_sc_hd__a22o_1 _24148_ (.A1(\decoded_imm_uj[5] ),
    .A2(_20031_),
    .B1(_20047_),
    .B2(\mem_rdata_q[25] ),
    .X(_20048_));
 sky130_fd_sc_hd__buf_2 _24149_ (.A(_18647_),
    .X(_20049_));
 sky130_fd_sc_hd__mux2_1 _24150_ (.A0(_20048_),
    .A1(\decoded_imm[5] ),
    .S(_20049_),
    .X(_02734_));
 sky130_fd_sc_hd__a22o_1 _24151_ (.A1(\decoded_imm_uj[6] ),
    .A2(_20031_),
    .B1(_20047_),
    .B2(_19737_),
    .X(_20050_));
 sky130_fd_sc_hd__mux2_1 _24152_ (.A0(_20050_),
    .A1(\decoded_imm[6] ),
    .S(_20049_),
    .X(_02733_));
 sky130_fd_sc_hd__a22o_1 _24153_ (.A1(\decoded_imm_uj[7] ),
    .A2(_20031_),
    .B1(_20047_),
    .B2(\mem_rdata_q[27] ),
    .X(_20051_));
 sky130_fd_sc_hd__mux2_1 _24154_ (.A0(_20051_),
    .A1(\decoded_imm[7] ),
    .S(_20049_),
    .X(_02732_));
 sky130_fd_sc_hd__a22o_1 _24155_ (.A1(\decoded_imm_uj[8] ),
    .A2(_20023_),
    .B1(_20047_),
    .B2(\mem_rdata_q[28] ),
    .X(_20052_));
 sky130_fd_sc_hd__mux2_1 _24156_ (.A0(_20052_),
    .A1(\decoded_imm[8] ),
    .S(_20049_),
    .X(_02731_));
 sky130_fd_sc_hd__a22o_1 _24157_ (.A1(\decoded_imm_uj[9] ),
    .A2(_20023_),
    .B1(_20047_),
    .B2(\mem_rdata_q[29] ),
    .X(_20053_));
 sky130_fd_sc_hd__mux2_1 _24158_ (.A0(_20053_),
    .A1(\decoded_imm[9] ),
    .S(_20049_),
    .X(_02730_));
 sky130_fd_sc_hd__a22o_1 _24159_ (.A1(\decoded_imm_uj[10] ),
    .A2(_20023_),
    .B1(_20047_),
    .B2(\mem_rdata_q[30] ),
    .X(_20054_));
 sky130_fd_sc_hd__mux2_1 _24160_ (.A0(_20054_),
    .A1(\decoded_imm[10] ),
    .S(_20049_),
    .X(_02729_));
 sky130_vsdinv _24161_ (.A(is_sb_sh_sw),
    .Y(_20055_));
 sky130_fd_sc_hd__a21oi_1 _24162_ (.A1(_19723_),
    .A2(_20055_),
    .B1(_18658_),
    .Y(_20056_));
 sky130_fd_sc_hd__a221o_2 _24163_ (.A1(is_beq_bne_blt_bge_bltu_bgeu),
    .A2(\mem_rdata_q[7] ),
    .B1(\decoded_imm_uj[11] ),
    .B2(_20022_),
    .C1(_20056_),
    .X(_20057_));
 sky130_fd_sc_hd__buf_2 _24164_ (.A(_18647_),
    .X(_20058_));
 sky130_fd_sc_hd__mux2_1 _24165_ (.A0(_20057_),
    .A1(\decoded_imm[11] ),
    .S(_20058_),
    .X(_02728_));
 sky130_vsdinv _24166_ (.A(_18503_),
    .Y(_20059_));
 sky130_fd_sc_hd__clkbuf_2 _24167_ (.A(_20059_),
    .X(_20060_));
 sky130_fd_sc_hd__and2_1 _24168_ (.A(_20046_),
    .B(_18672_),
    .X(_20061_));
 sky130_fd_sc_hd__buf_2 _24169_ (.A(_20061_),
    .X(_20062_));
 sky130_fd_sc_hd__a221o_2 _24170_ (.A1(\decoded_imm_uj[12] ),
    .A2(_20023_),
    .B1(_18692_),
    .B2(_20060_),
    .C1(_20062_),
    .X(_20063_));
 sky130_fd_sc_hd__mux2_1 _24171_ (.A0(_20063_),
    .A1(\decoded_imm[12] ),
    .S(_20058_),
    .X(_02727_));
 sky130_fd_sc_hd__buf_2 _24172_ (.A(_20022_),
    .X(_20064_));
 sky130_fd_sc_hd__a221o_2 _24173_ (.A1(\decoded_imm_uj[13] ),
    .A2(_20064_),
    .B1(\mem_rdata_q[13] ),
    .B2(_20060_),
    .C1(_20062_),
    .X(_20065_));
 sky130_fd_sc_hd__mux2_1 _24174_ (.A0(_20065_),
    .A1(\decoded_imm[13] ),
    .S(_20058_),
    .X(_02726_));
 sky130_fd_sc_hd__buf_2 _24175_ (.A(_20059_),
    .X(_20066_));
 sky130_fd_sc_hd__a221o_1 _24176_ (.A1(\decoded_imm_uj[14] ),
    .A2(_20064_),
    .B1(_18667_),
    .B2(_20066_),
    .C1(_20062_),
    .X(_20067_));
 sky130_fd_sc_hd__mux2_1 _24177_ (.A0(_20067_),
    .A1(\decoded_imm[14] ),
    .S(_20058_),
    .X(_02725_));
 sky130_fd_sc_hd__a221o_1 _24178_ (.A1(\decoded_imm_uj[15] ),
    .A2(_20064_),
    .B1(\mem_rdata_q[15] ),
    .B2(_20066_),
    .C1(_20062_),
    .X(_20068_));
 sky130_fd_sc_hd__mux2_1 _24179_ (.A0(_20068_),
    .A1(\decoded_imm[15] ),
    .S(_20058_),
    .X(_02724_));
 sky130_fd_sc_hd__a221o_1 _24180_ (.A1(\decoded_imm_uj[16] ),
    .A2(_20064_),
    .B1(\mem_rdata_q[16] ),
    .B2(_20066_),
    .C1(_20062_),
    .X(_20069_));
 sky130_fd_sc_hd__mux2_1 _24181_ (.A0(_20069_),
    .A1(\decoded_imm[16] ),
    .S(_20058_),
    .X(_02723_));
 sky130_fd_sc_hd__a221o_1 _24182_ (.A1(\decoded_imm_uj[17] ),
    .A2(_20064_),
    .B1(\mem_rdata_q[17] ),
    .B2(_20066_),
    .C1(_20062_),
    .X(_20070_));
 sky130_fd_sc_hd__mux2_1 _24183_ (.A0(_20070_),
    .A1(\decoded_imm[17] ),
    .S(_20034_),
    .X(_02722_));
 sky130_fd_sc_hd__a221o_1 _24184_ (.A1(\decoded_imm_uj[18] ),
    .A2(_20064_),
    .B1(\mem_rdata_q[18] ),
    .B2(_20066_),
    .C1(_20061_),
    .X(_20071_));
 sky130_fd_sc_hd__mux2_1 _24185_ (.A0(_20071_),
    .A1(\decoded_imm[18] ),
    .S(_20034_),
    .X(_02721_));
 sky130_fd_sc_hd__a221o_1 _24186_ (.A1(\decoded_imm_uj[19] ),
    .A2(_20022_),
    .B1(\mem_rdata_q[19] ),
    .B2(_20066_),
    .C1(_20061_),
    .X(_20072_));
 sky130_fd_sc_hd__mux2_1 _24187_ (.A0(_20072_),
    .A1(\decoded_imm[19] ),
    .S(_20034_),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_2 _24188_ (.A(_18503_),
    .X(_20073_));
 sky130_fd_sc_hd__buf_1 _24189_ (.A(_19700_),
    .X(_20074_));
 sky130_fd_sc_hd__o21ai_1 _24190_ (.A1(_19720_),
    .A2(_20073_),
    .B1(_20074_),
    .Y(_20075_));
 sky130_fd_sc_hd__nor2_2 _24191_ (.A(_18658_),
    .B(_19723_),
    .Y(_20076_));
 sky130_fd_sc_hd__clkbuf_2 _24192_ (.A(_20076_),
    .X(_20077_));
 sky130_vsdinv _24193_ (.A(\decoded_imm_uj[20] ),
    .Y(_20078_));
 sky130_fd_sc_hd__clkbuf_4 _24194_ (.A(_20078_),
    .X(_20079_));
 sky130_fd_sc_hd__buf_4 _24195_ (.A(_20079_),
    .X(_20080_));
 sky130_fd_sc_hd__o22a_1 _24196_ (.A1(_20080_),
    .A2(_00323_),
    .B1(_18658_),
    .B2(_20025_),
    .X(_20081_));
 sky130_vsdinv _24197_ (.A(_20081_),
    .Y(_20082_));
 sky130_fd_sc_hd__clkbuf_2 _24198_ (.A(_20082_),
    .X(_20083_));
 sky130_fd_sc_hd__o32a_1 _24199_ (.A1(_20075_),
    .A2(_20077_),
    .A3(_20083_),
    .B1(\decoded_imm[20] ),
    .B2(_19777_),
    .X(_02719_));
 sky130_fd_sc_hd__o21ai_1 _24200_ (.A1(_19764_),
    .A2(_20073_),
    .B1(_20074_),
    .Y(_20084_));
 sky130_fd_sc_hd__nor2_1 _24201_ (.A(_20076_),
    .B(_20082_),
    .Y(_20085_));
 sky130_vsdinv _24202_ (.A(_20085_),
    .Y(_20086_));
 sky130_fd_sc_hd__o22a_1 _24203_ (.A1(\decoded_imm[21] ),
    .A2(_19699_),
    .B1(_20084_),
    .B2(_20086_),
    .X(_02718_));
 sky130_fd_sc_hd__a21o_1 _24204_ (.A1(\mem_rdata_q[22] ),
    .A2(_20060_),
    .B1(_18711_),
    .X(_20087_));
 sky130_fd_sc_hd__o32a_1 _24205_ (.A1(_20083_),
    .A2(_20077_),
    .A3(_20087_),
    .B1(\decoded_imm[22] ),
    .B2(_19777_),
    .X(_02717_));
 sky130_fd_sc_hd__a21o_1 _24206_ (.A1(\mem_rdata_q[23] ),
    .A2(_20060_),
    .B1(_18711_),
    .X(_20088_));
 sky130_fd_sc_hd__clkbuf_2 _24207_ (.A(_18728_),
    .X(_20089_));
 sky130_fd_sc_hd__o32a_1 _24208_ (.A1(_20083_),
    .A2(_20077_),
    .A3(_20088_),
    .B1(\decoded_imm[23] ),
    .B2(_20089_),
    .X(_02716_));
 sky130_fd_sc_hd__a21o_1 _24209_ (.A1(\mem_rdata_q[24] ),
    .A2(_20060_),
    .B1(_18647_),
    .X(_20090_));
 sky130_fd_sc_hd__o32a_1 _24210_ (.A1(_20083_),
    .A2(_20077_),
    .A3(_20090_),
    .B1(\decoded_imm[24] ),
    .B2(_20089_),
    .X(_02715_));
 sky130_fd_sc_hd__o21ai_1 _24211_ (.A1(_18656_),
    .A2(_20073_),
    .B1(_20074_),
    .Y(_20091_));
 sky130_fd_sc_hd__o32a_1 _24212_ (.A1(_20091_),
    .A2(_20077_),
    .A3(_20083_),
    .B1(\decoded_imm[25] ),
    .B2(_20089_),
    .X(_02714_));
 sky130_fd_sc_hd__a21o_1 _24213_ (.A1(_19737_),
    .A2(_20060_),
    .B1(_18690_),
    .X(_20092_));
 sky130_fd_sc_hd__o22a_1 _24214_ (.A1(\decoded_imm[26] ),
    .A2(_19699_),
    .B1(_20092_),
    .B2(_20086_),
    .X(_02713_));
 sky130_fd_sc_hd__o21ai_1 _24215_ (.A1(_18655_),
    .A2(_20073_),
    .B1(_20074_),
    .Y(_20093_));
 sky130_fd_sc_hd__o32a_1 _24216_ (.A1(_20093_),
    .A2(_20077_),
    .A3(_20083_),
    .B1(\decoded_imm[27] ),
    .B2(_20089_),
    .X(_02712_));
 sky130_fd_sc_hd__o21ai_1 _24217_ (.A1(_19736_),
    .A2(_20073_),
    .B1(_20074_),
    .Y(_20094_));
 sky130_fd_sc_hd__o32a_1 _24218_ (.A1(_20094_),
    .A2(_20076_),
    .A3(_20082_),
    .B1(\decoded_imm[28] ),
    .B2(_20089_),
    .X(_02711_));
 sky130_fd_sc_hd__o21ai_1 _24219_ (.A1(_18660_),
    .A2(_20073_),
    .B1(_20074_),
    .Y(_20095_));
 sky130_fd_sc_hd__o22a_1 _24220_ (.A1(\decoded_imm[29] ),
    .A2(_19701_),
    .B1(_20095_),
    .B2(_20086_),
    .X(_02710_));
 sky130_fd_sc_hd__o21ai_1 _24221_ (.A1(_18659_),
    .A2(_18503_),
    .B1(_18728_),
    .Y(_20096_));
 sky130_fd_sc_hd__o32a_1 _24222_ (.A1(_20096_),
    .A2(_20076_),
    .A3(_20082_),
    .B1(\decoded_imm[30] ),
    .B2(_20089_),
    .X(_02709_));
 sky130_fd_sc_hd__or2_1 _24223_ (.A(_20059_),
    .B(_20046_),
    .X(_20097_));
 sky130_fd_sc_hd__a22o_1 _24224_ (.A1(_19711_),
    .A2(_20023_),
    .B1(_20097_),
    .B2(_18672_),
    .X(_20098_));
 sky130_fd_sc_hd__mux2_1 _24225_ (.A0(_20098_),
    .A1(\decoded_imm[31] ),
    .S(_20034_),
    .X(_02708_));
 sky130_fd_sc_hd__and3_4 _24226_ (.A(_19489_),
    .B(_18542_),
    .C(_19488_),
    .X(_20099_));
 sky130_fd_sc_hd__clkbuf_2 _24227_ (.A(_20099_),
    .X(_20100_));
 sky130_fd_sc_hd__nor2_1 _24228_ (.A(_19365_),
    .B(_20100_),
    .Y(_20101_));
 sky130_fd_sc_hd__a31o_1 _24229_ (.A1(_20890_),
    .A2(_18539_),
    .A3(_20100_),
    .B1(_20101_),
    .X(_02707_));
 sky130_fd_sc_hd__buf_6 _24230_ (.A(_18446_),
    .X(_00308_));
 sky130_fd_sc_hd__nor2_8 _24231_ (.A(_02542_),
    .B(_00308_),
    .Y(_20102_));
 sky130_fd_sc_hd__nor2_1 _24232_ (.A(_19364_),
    .B(_20100_),
    .Y(_20103_));
 sky130_fd_sc_hd__a31o_1 _24233_ (.A1(_20102_),
    .A2(\decoded_rd[1] ),
    .A3(_20100_),
    .B1(_20103_),
    .X(_02706_));
 sky130_fd_sc_hd__nor2_1 _24234_ (.A(_19463_),
    .B(_20099_),
    .Y(_20104_));
 sky130_fd_sc_hd__a31o_1 _24235_ (.A1(_20102_),
    .A2(\decoded_rd[2] ),
    .A3(_20100_),
    .B1(_20104_),
    .X(_02705_));
 sky130_fd_sc_hd__nor2_1 _24236_ (.A(_19368_),
    .B(_20099_),
    .Y(_20105_));
 sky130_fd_sc_hd__a31o_1 _24237_ (.A1(_20102_),
    .A2(\decoded_rd[3] ),
    .A3(_20100_),
    .B1(_20105_),
    .X(_02704_));
 sky130_fd_sc_hd__or3_1 _24238_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(is_slli_srli_srai),
    .C(is_lui_auipc_jal),
    .X(_20106_));
 sky130_vsdinv _24239_ (.A(_20106_),
    .Y(_20107_));
 sky130_fd_sc_hd__nor2_1 _24240_ (.A(_18543_),
    .B(_20107_),
    .Y(_20108_));
 sky130_fd_sc_hd__and3_1 _24241_ (.A(_18547_),
    .B(_20055_),
    .C(_18519_),
    .X(_20109_));
 sky130_fd_sc_hd__o21a_1 _24242_ (.A1(_20108_),
    .A2(_20109_),
    .B1(_19427_),
    .X(_02703_));
 sky130_vsdinv _24243_ (.A(net226),
    .Y(_20110_));
 sky130_fd_sc_hd__clkbuf_2 _24244_ (.A(_20110_),
    .X(_20111_));
 sky130_fd_sc_hd__buf_2 _24245_ (.A(_20111_),
    .X(_02327_));
 sky130_fd_sc_hd__and2_1 _24246_ (.A(_02327_),
    .B(_02558_),
    .X(_02702_));
 sky130_fd_sc_hd__and2_1 _24247_ (.A(_02327_),
    .B(_02557_),
    .X(_02701_));
 sky130_fd_sc_hd__and2_1 _24248_ (.A(_02327_),
    .B(_02556_),
    .X(_02700_));
 sky130_fd_sc_hd__and2_1 _24249_ (.A(_02327_),
    .B(_02555_),
    .X(_02699_));
 sky130_fd_sc_hd__and2_1 _24250_ (.A(_20111_),
    .B(_02554_),
    .X(_02698_));
 sky130_fd_sc_hd__and2_1 _24251_ (.A(_20111_),
    .B(_02553_),
    .X(_02697_));
 sky130_fd_sc_hd__and2_1 _24252_ (.A(_20111_),
    .B(_02552_),
    .X(_02696_));
 sky130_fd_sc_hd__and2_1 _24253_ (.A(_20111_),
    .B(_02551_),
    .X(_02695_));
 sky130_vsdinv _24254_ (.A(net225),
    .Y(_20112_));
 sky130_fd_sc_hd__clkbuf_2 _24255_ (.A(_20112_),
    .X(_02324_));
 sky130_fd_sc_hd__and2_1 _24256_ (.A(_02324_),
    .B(_00122_),
    .X(_02550_));
 sky130_fd_sc_hd__nor2_1 _24257_ (.A(net226),
    .B(net225),
    .Y(_20113_));
 sky130_fd_sc_hd__buf_1 _24258_ (.A(_20113_),
    .X(_20114_));
 sky130_fd_sc_hd__and2_1 _24259_ (.A(_20114_),
    .B(_00122_),
    .X(_02694_));
 sky130_fd_sc_hd__and2_1 _24260_ (.A(_02324_),
    .B(_00116_),
    .X(_02549_));
 sky130_fd_sc_hd__and2_1 _24261_ (.A(_20114_),
    .B(_00116_),
    .X(_02693_));
 sky130_fd_sc_hd__and2_1 _24262_ (.A(_02324_),
    .B(_00110_),
    .X(_02548_));
 sky130_fd_sc_hd__and2_1 _24263_ (.A(_20114_),
    .B(_00110_),
    .X(_02692_));
 sky130_fd_sc_hd__and2_1 _24264_ (.A(_02324_),
    .B(_00104_),
    .X(_02547_));
 sky130_fd_sc_hd__and2_1 _24265_ (.A(_20114_),
    .B(_00104_),
    .X(_02691_));
 sky130_fd_sc_hd__nor2_2 _24266_ (.A(_19451_),
    .B(_19452_),
    .Y(_20115_));
 sky130_fd_sc_hd__and2_1 _24267_ (.A(_20115_),
    .B(_00094_),
    .X(_02546_));
 sky130_vsdinv _24268_ (.A(net222),
    .Y(_20116_));
 sky130_fd_sc_hd__buf_2 _24269_ (.A(_20116_),
    .X(_02321_));
 sky130_fd_sc_hd__and3_1 _24270_ (.A(_20114_),
    .B(_02321_),
    .C(_00094_),
    .X(_02690_));
 sky130_fd_sc_hd__and2_1 _24271_ (.A(_20115_),
    .B(_00084_),
    .X(_02545_));
 sky130_fd_sc_hd__and3_1 _24272_ (.A(_20113_),
    .B(_02321_),
    .C(_00084_),
    .X(_02689_));
 sky130_vsdinv _24273_ (.A(net211),
    .Y(_20117_));
 sky130_fd_sc_hd__buf_2 _24274_ (.A(_20117_),
    .X(_02318_));
 sky130_fd_sc_hd__and3_1 _24275_ (.A(_20115_),
    .B(_02318_),
    .C(_00066_),
    .X(_02544_));
 sky130_fd_sc_hd__and3_1 _24276_ (.A(_20116_),
    .B(_02318_),
    .C(_00066_),
    .X(_00068_));
 sky130_fd_sc_hd__and2_1 _24277_ (.A(_00068_),
    .B(_20114_),
    .X(_02688_));
 sky130_vsdinv _24278_ (.A(net306),
    .Y(_20118_));
 sky130_fd_sc_hd__buf_4 _24279_ (.A(_20118_),
    .X(_20119_));
 sky130_fd_sc_hd__nor2_1 _24280_ (.A(net211),
    .B(net200),
    .Y(_20120_));
 sky130_fd_sc_hd__and2_1 _24281_ (.A(_20120_),
    .B(_20116_),
    .X(_20121_));
 sky130_fd_sc_hd__nand2_1 _24282_ (.A(_20121_),
    .B(_20112_),
    .Y(_20122_));
 sky130_fd_sc_hd__nor2_1 _24283_ (.A(_20119_),
    .B(_20122_),
    .Y(_02543_));
 sky130_fd_sc_hd__and2_1 _24284_ (.A(_02543_),
    .B(_20111_),
    .X(_02687_));
 sky130_fd_sc_hd__o211a_1 _24285_ (.A1(\reg_pc[1] ),
    .A2(\reg_next_pc[0] ),
    .B1(net101),
    .C1(_18346_),
    .X(_20123_));
 sky130_fd_sc_hd__clkbuf_4 _24286_ (.A(_20123_),
    .X(_00307_));
 sky130_fd_sc_hd__and3_1 _24287_ (.A(_18449_),
    .B(_18579_),
    .C(_18623_),
    .X(_00312_));
 sky130_fd_sc_hd__nor2_2 _24288_ (.A(_18308_),
    .B(_18319_),
    .Y(_00303_));
 sky130_vsdinv _24289_ (.A(_00303_),
    .Y(_20124_));
 sky130_fd_sc_hd__nor2_1 _24290_ (.A(_00307_),
    .B(_20124_),
    .Y(_20125_));
 sky130_vsdinv _24291_ (.A(_00308_),
    .Y(_20126_));
 sky130_fd_sc_hd__or2_1 _24292_ (.A(instr_waitirq),
    .B(_18381_),
    .X(_20127_));
 sky130_fd_sc_hd__nand2_2 _24293_ (.A(_18449_),
    .B(_18625_),
    .Y(_20128_));
 sky130_fd_sc_hd__nor3_4 _24294_ (.A(\pcpi_mul.active[1] ),
    .B(_00311_),
    .C(_20128_),
    .Y(_20129_));
 sky130_fd_sc_hd__nor2_1 _24295_ (.A(_18311_),
    .B(_19147_),
    .Y(_20130_));
 sky130_fd_sc_hd__a32o_1 _24296_ (.A1(_20126_),
    .A2(_19370_),
    .A3(_20127_),
    .B1(_20129_),
    .B2(_20130_),
    .X(_20131_));
 sky130_vsdinv _24297_ (.A(\mem_wordsize[2] ),
    .Y(_20132_));
 sky130_fd_sc_hd__nor2_4 _24298_ (.A(_20118_),
    .B(_20132_),
    .Y(_00306_));
 sky130_fd_sc_hd__nor2_2 _24299_ (.A(irq_active),
    .B(\irq_mask[2] ),
    .Y(_20133_));
 sky130_fd_sc_hd__clkbuf_2 _24300_ (.A(_20133_),
    .X(_20134_));
 sky130_vsdinv _24301_ (.A(\mem_wordsize[0] ),
    .Y(_20135_));
 sky130_fd_sc_hd__nor2_8 _24302_ (.A(_19818_),
    .B(_19820_),
    .Y(_00304_));
 sky130_fd_sc_hd__nor2_8 _24303_ (.A(_20135_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__nor2_2 _24304_ (.A(_00306_),
    .B(_00305_),
    .Y(_20136_));
 sky130_fd_sc_hd__or2_1 _24305_ (.A(_20134_),
    .B(_20136_),
    .X(_20137_));
 sky130_fd_sc_hd__a32o_1 _24306_ (.A1(_20131_),
    .A2(_00306_),
    .A3(_20134_),
    .B1(_03828_),
    .B2(_20137_),
    .X(_20138_));
 sky130_vsdinv _24307_ (.A(_20123_),
    .Y(_20139_));
 sky130_fd_sc_hd__o21a_1 _24308_ (.A1(_20124_),
    .A2(_20136_),
    .B1(_20139_),
    .X(_20140_));
 sky130_fd_sc_hd__nor2_4 _24309_ (.A(_20134_),
    .B(_20140_),
    .Y(_20141_));
 sky130_vsdinv _24310_ (.A(_20133_),
    .Y(_20142_));
 sky130_fd_sc_hd__nor2_1 _24311_ (.A(_20142_),
    .B(_00306_),
    .Y(_20143_));
 sky130_vsdinv _24312_ (.A(_00305_),
    .Y(_20144_));
 sky130_fd_sc_hd__nor2_1 _24313_ (.A(_20144_),
    .B(_20124_),
    .Y(_20145_));
 sky130_fd_sc_hd__nor2_2 _24314_ (.A(_20142_),
    .B(_20139_),
    .Y(_20146_));
 sky130_fd_sc_hd__or2_1 _24315_ (.A(_20146_),
    .B(_20140_),
    .X(_20147_));
 sky130_fd_sc_hd__a31o_1 _24316_ (.A1(_20139_),
    .A2(_20143_),
    .A3(_20145_),
    .B1(_20147_),
    .X(_20148_));
 sky130_fd_sc_hd__a2bb2o_1 _24317_ (.A1_N(_18462_),
    .A2_N(_20141_),
    .B1(_20129_),
    .B2(_20148_),
    .X(_20149_));
 sky130_fd_sc_hd__buf_2 _24318_ (.A(_18519_),
    .X(_20150_));
 sky130_fd_sc_hd__and3_1 _24319_ (.A(_00310_),
    .B(_20149_),
    .C(_20150_),
    .X(_20151_));
 sky130_fd_sc_hd__a22o_1 _24320_ (.A1(_00309_),
    .A2(_20146_),
    .B1(_00308_),
    .B2(_20147_),
    .X(_20152_));
 sky130_fd_sc_hd__nor2_1 _24321_ (.A(_18542_),
    .B(_18495_),
    .Y(_20153_));
 sky130_fd_sc_hd__o21a_1 _24322_ (.A1(_18481_),
    .A2(_18323_),
    .B1(_18540_),
    .X(_20154_));
 sky130_fd_sc_hd__o21a_1 _24323_ (.A1(_18319_),
    .A2(_00307_),
    .B1(_03828_),
    .X(_20155_));
 sky130_fd_sc_hd__nor2_2 _24324_ (.A(_18319_),
    .B(_20136_),
    .Y(_20156_));
 sky130_fd_sc_hd__o21ai_2 _24325_ (.A1(_00307_),
    .A2(_20156_),
    .B1(_20142_),
    .Y(_20157_));
 sky130_fd_sc_hd__o31a_1 _24326_ (.A1(_20153_),
    .A2(_20154_),
    .A3(_20155_),
    .B1(_20157_),
    .X(_20158_));
 sky130_fd_sc_hd__a2111o_1 _24327_ (.A1(_20152_),
    .A2(_18754_),
    .B1(_18578_),
    .C1(_00314_),
    .D1(_20158_),
    .X(_20159_));
 sky130_fd_sc_hd__and3_1 _24328_ (.A(_18447_),
    .B(_20022_),
    .C(decoder_trigger),
    .X(_20160_));
 sky130_fd_sc_hd__clkbuf_1 _24329_ (.A(_20160_),
    .X(_02062_));
 sky130_fd_sc_hd__nand2_1 _24330_ (.A(_02062_),
    .B(_18330_),
    .Y(_20161_));
 sky130_vsdinv _24331_ (.A(_00306_),
    .Y(_20162_));
 sky130_fd_sc_hd__nand2_1 _24332_ (.A(_00303_),
    .B(_20133_),
    .Y(_20163_));
 sky130_fd_sc_hd__o22a_1 _24333_ (.A1(_20142_),
    .A2(_20139_),
    .B1(_20162_),
    .B2(_20163_),
    .X(_20164_));
 sky130_fd_sc_hd__and3_1 _24334_ (.A(_19163_),
    .B(_18381_),
    .C(_19162_),
    .X(_20165_));
 sky130_fd_sc_hd__nand2_1 _24335_ (.A(_20165_),
    .B(_20146_),
    .Y(_20166_));
 sky130_fd_sc_hd__nand2_1 _24336_ (.A(_20125_),
    .B(_20162_),
    .Y(_20167_));
 sky130_fd_sc_hd__a2111o_1 _24337_ (.A1(_20142_),
    .A2(_00305_),
    .B1(_19162_),
    .C1(_20167_),
    .D1(_19164_),
    .X(_20168_));
 sky130_vsdinv _24338_ (.A(_20143_),
    .Y(_20169_));
 sky130_fd_sc_hd__o32a_1 _24339_ (.A1(_20126_),
    .A2(_20136_),
    .A3(_20163_),
    .B1(_20169_),
    .B2(_20161_),
    .X(_20170_));
 sky130_fd_sc_hd__o32a_1 _24340_ (.A1(_19162_),
    .A2(_19164_),
    .A3(_00303_),
    .B1(_20156_),
    .B2(_20161_),
    .X(_20171_));
 sky130_vsdinv _24341_ (.A(_20156_),
    .Y(_20172_));
 sky130_vsdinv _24342_ (.A(_20145_),
    .Y(_20173_));
 sky130_fd_sc_hd__nor2_1 _24343_ (.A(_20169_),
    .B(_20173_),
    .Y(_20174_));
 sky130_fd_sc_hd__o21ai_1 _24344_ (.A1(_20172_),
    .A2(_20174_),
    .B1(_20165_),
    .Y(_20175_));
 sky130_fd_sc_hd__a31o_1 _24345_ (.A1(_20170_),
    .A2(_20171_),
    .A3(_20175_),
    .B1(_00307_),
    .X(_20176_));
 sky130_fd_sc_hd__o2111a_1 _24346_ (.A1(_20161_),
    .A2(_20164_),
    .B1(_20166_),
    .C1(_20168_),
    .D1(_20176_),
    .X(_20177_));
 sky130_fd_sc_hd__nor2_1 _24347_ (.A(_18528_),
    .B(_20177_),
    .Y(_20178_));
 sky130_fd_sc_hd__a2111o_1 _24348_ (.A1(_20125_),
    .A2(_20138_),
    .B1(_20151_),
    .C1(_20159_),
    .D1(_20178_),
    .X(_00039_));
 sky130_fd_sc_hd__nor2_1 _24349_ (.A(_18532_),
    .B(_20141_),
    .Y(_20179_));
 sky130_vsdinv _24350_ (.A(_20179_),
    .Y(_20180_));
 sky130_fd_sc_hd__nor2_1 _24351_ (.A(_20180_),
    .B(_18560_),
    .Y(_00040_));
 sky130_fd_sc_hd__nand2_1 _24352_ (.A(_18545_),
    .B(_18496_),
    .Y(_20181_));
 sky130_fd_sc_hd__clkbuf_2 _24353_ (.A(_18328_),
    .X(_20182_));
 sky130_fd_sc_hd__clkbuf_4 _24354_ (.A(_20182_),
    .X(_20183_));
 sky130_fd_sc_hd__or2_1 _24355_ (.A(_20183_),
    .B(_19167_),
    .X(_20184_));
 sky130_fd_sc_hd__a21oi_1 _24356_ (.A1(_20181_),
    .A2(_20184_),
    .B1(_20180_),
    .Y(_00044_));
 sky130_fd_sc_hd__a32o_1 _24357_ (.A1(_18546_),
    .A2(_18495_),
    .A3(_20107_),
    .B1(_19145_),
    .B2(_19146_),
    .X(_20185_));
 sky130_fd_sc_hd__and2_1 _24358_ (.A(_20185_),
    .B(_20179_),
    .X(_00041_));
 sky130_fd_sc_hd__or4b_4 _24359_ (.A(\pcpi_mul.active[1] ),
    .B(_00311_),
    .C(_19147_),
    .D_N(_20128_),
    .X(_20186_));
 sky130_fd_sc_hd__a31oi_1 _24360_ (.A1(_20186_),
    .A2(_19362_),
    .A3(_20157_),
    .B1(_18870_),
    .Y(_00038_));
 sky130_fd_sc_hd__nor2_1 _24361_ (.A(_18312_),
    .B(_18557_),
    .Y(_20187_));
 sky130_vsdinv _24362_ (.A(_20187_),
    .Y(_20188_));
 sky130_fd_sc_hd__or3_1 _24363_ (.A(_18311_),
    .B(_20055_),
    .C(_18520_),
    .X(_20189_));
 sky130_fd_sc_hd__o32a_1 _24364_ (.A1(_19782_),
    .A2(_20173_),
    .A3(_20188_),
    .B1(_20163_),
    .B2(_20189_),
    .X(_20190_));
 sky130_fd_sc_hd__nor2_1 _24365_ (.A(_20144_),
    .B(_20167_),
    .Y(_20191_));
 sky130_fd_sc_hd__o32a_1 _24366_ (.A1(_18311_),
    .A2(_18324_),
    .A3(_19167_),
    .B1(_20191_),
    .B2(_20188_),
    .X(_20192_));
 sky130_fd_sc_hd__o22a_1 _24367_ (.A1(_20191_),
    .A2(_20189_),
    .B1(_19782_),
    .B2(_20192_),
    .X(_20193_));
 sky130_fd_sc_hd__o32ai_4 _24368_ (.A1(_00307_),
    .A2(_20169_),
    .A3(_20190_),
    .B1(_20141_),
    .B2(_20193_),
    .Y(_00043_));
 sky130_fd_sc_hd__o21a_4 _24369_ (.A1(mem_do_rdata),
    .A2(_18348_),
    .B1(_19472_),
    .X(net199));
 sky130_fd_sc_hd__nand2_2 _24370_ (.A(_18350_),
    .B(_19472_),
    .Y(_00316_));
 sky130_fd_sc_hd__nor2_1 _24371_ (.A(_00291_),
    .B(_19782_),
    .Y(_00317_));
 sky130_fd_sc_hd__clkbuf_4 _24372_ (.A(_18487_),
    .X(_20194_));
 sky130_fd_sc_hd__buf_2 _24373_ (.A(_20194_),
    .X(_20195_));
 sky130_fd_sc_hd__o21a_1 _24374_ (.A1(_00305_),
    .A2(_20167_),
    .B1(_20164_),
    .X(_20196_));
 sky130_fd_sc_hd__o32a_1 _24375_ (.A1(_18554_),
    .A2(_20196_),
    .A3(_18557_),
    .B1(_00302_),
    .B2(_20180_),
    .X(_20197_));
 sky130_fd_sc_hd__or2_1 _24376_ (.A(_20124_),
    .B(_20174_),
    .X(_20198_));
 sky130_fd_sc_hd__and3_1 _24377_ (.A(_20139_),
    .B(\cpu_state[4] ),
    .C(_18482_),
    .X(_20199_));
 sky130_fd_sc_hd__o21a_1 _24378_ (.A1(_20108_),
    .A2(_20109_),
    .B1(_20157_),
    .X(_20200_));
 sky130_fd_sc_hd__a31o_1 _24379_ (.A1(_18322_),
    .A2(_20198_),
    .A3(_20199_),
    .B1(_20200_),
    .X(_20201_));
 sky130_fd_sc_hd__a2bb2o_1 _24380_ (.A1_N(_20195_),
    .A2_N(_20197_),
    .B1(_18696_),
    .B2(_20201_),
    .X(_00042_));
 sky130_fd_sc_hd__nor2_2 _24381_ (.A(net200),
    .B(_20118_),
    .Y(_00048_));
 sky130_vsdinv _24382_ (.A(net200),
    .Y(_20202_));
 sky130_fd_sc_hd__nor2_2 _24383_ (.A(net306),
    .B(_20202_),
    .Y(_20203_));
 sky130_fd_sc_hd__or2_2 _24384_ (.A(_00048_),
    .B(_20203_),
    .X(_02591_));
 sky130_fd_sc_hd__nor2_1 _24385_ (.A(net355),
    .B(net323),
    .Y(_20204_));
 sky130_fd_sc_hd__inv_2 _24386_ (.A(net355),
    .Y(_02390_));
 sky130_vsdinv _24387_ (.A(net323),
    .Y(_20205_));
 sky130_fd_sc_hd__nor2_2 _24388_ (.A(_02390_),
    .B(_20205_),
    .Y(_20206_));
 sky130_fd_sc_hd__nor2_1 _24389_ (.A(_20204_),
    .B(_20206_),
    .Y(_20207_));
 sky130_vsdinv _24390_ (.A(_20207_),
    .Y(_20208_));
 sky130_fd_sc_hd__nor2_1 _24391_ (.A(net356),
    .B(net324),
    .Y(_20209_));
 sky130_fd_sc_hd__inv_2 _24392_ (.A(net356),
    .Y(_02393_));
 sky130_vsdinv _24393_ (.A(net324),
    .Y(_20210_));
 sky130_fd_sc_hd__nor2_2 _24394_ (.A(_02393_),
    .B(_20210_),
    .Y(_20211_));
 sky130_fd_sc_hd__or2_1 _24395_ (.A(_20209_),
    .B(_20211_),
    .X(_20212_));
 sky130_fd_sc_hd__nor2_1 _24396_ (.A(net357),
    .B(net325),
    .Y(_20213_));
 sky130_vsdinv _24397_ (.A(_20213_),
    .Y(_20214_));
 sky130_fd_sc_hd__nand2_1 _24398_ (.A(_19429_),
    .B(net325),
    .Y(_20215_));
 sky130_fd_sc_hd__nand2_1 _24399_ (.A(_20214_),
    .B(_20215_),
    .Y(_20216_));
 sky130_fd_sc_hd__inv_2 _24400_ (.A(net354),
    .Y(_02387_));
 sky130_vsdinv _24401_ (.A(net322),
    .Y(_20217_));
 sky130_fd_sc_hd__nand2_1 _24402_ (.A(_02387_),
    .B(_20217_),
    .Y(_20218_));
 sky130_fd_sc_hd__nand2_1 _24403_ (.A(net354),
    .B(_19792_),
    .Y(_20219_));
 sky130_fd_sc_hd__nand2_1 _24404_ (.A(_20218_),
    .B(_20219_),
    .Y(_20220_));
 sky130_fd_sc_hd__and4_1 _24405_ (.A(_20208_),
    .B(_20212_),
    .C(_20216_),
    .D(_20220_),
    .X(_20221_));
 sky130_fd_sc_hd__nor2_1 _24406_ (.A(net330),
    .B(net362),
    .Y(_20222_));
 sky130_fd_sc_hd__nand2_1 _24407_ (.A(net330),
    .B(net362),
    .Y(_20223_));
 sky130_fd_sc_hd__or2b_2 _24408_ (.A(_20222_),
    .B_N(_20223_),
    .X(_20224_));
 sky130_fd_sc_hd__inv_2 _24409_ (.A(net361),
    .Y(_02405_));
 sky130_vsdinv _24410_ (.A(net329),
    .Y(_20225_));
 sky130_fd_sc_hd__nand2_1 _24411_ (.A(_02405_),
    .B(_20225_),
    .Y(_20226_));
 sky130_fd_sc_hd__nand2_1 _24412_ (.A(_19428_),
    .B(net329),
    .Y(_20227_));
 sky130_fd_sc_hd__nand2_1 _24413_ (.A(_20226_),
    .B(_20227_),
    .Y(_20228_));
 sky130_fd_sc_hd__and2_1 _24414_ (.A(_20224_),
    .B(_20228_),
    .X(_20229_));
 sky130_fd_sc_hd__nor2_1 _24415_ (.A(net359),
    .B(net327),
    .Y(_20230_));
 sky130_fd_sc_hd__inv_2 _24416_ (.A(net359),
    .Y(_02402_));
 sky130_vsdinv _24417_ (.A(net327),
    .Y(_20231_));
 sky130_fd_sc_hd__nor2_2 _24418_ (.A(_02402_),
    .B(_20231_),
    .Y(_20232_));
 sky130_fd_sc_hd__nor2_1 _24419_ (.A(_20230_),
    .B(_20232_),
    .Y(_20233_));
 sky130_vsdinv _24420_ (.A(_20233_),
    .Y(_20234_));
 sky130_fd_sc_hd__nor2_1 _24421_ (.A(net358),
    .B(net326),
    .Y(_20235_));
 sky130_fd_sc_hd__inv_2 _24422_ (.A(net358),
    .Y(_02399_));
 sky130_vsdinv _24423_ (.A(net326),
    .Y(_20236_));
 sky130_fd_sc_hd__nor2_2 _24424_ (.A(_02399_),
    .B(_20236_),
    .Y(_20237_));
 sky130_fd_sc_hd__nor2_1 _24425_ (.A(_20235_),
    .B(_20237_),
    .Y(_20238_));
 sky130_vsdinv _24426_ (.A(_20238_),
    .Y(_20239_));
 sky130_fd_sc_hd__and4_1 _24427_ (.A(_20221_),
    .B(_20229_),
    .C(_20234_),
    .D(_20239_),
    .X(_20240_));
 sky130_fd_sc_hd__nor2_1 _24428_ (.A(_19432_),
    .B(_19794_),
    .Y(_20241_));
 sky130_fd_sc_hd__inv_2 _24429_ (.A(net352),
    .Y(_02381_));
 sky130_vsdinv _24430_ (.A(net320),
    .Y(_20242_));
 sky130_fd_sc_hd__nor2_1 _24431_ (.A(_02381_),
    .B(_20242_),
    .Y(_20243_));
 sky130_fd_sc_hd__inv_2 _24432_ (.A(net350),
    .Y(_02375_));
 sky130_vsdinv _24433_ (.A(net318),
    .Y(_20244_));
 sky130_fd_sc_hd__nand2_1 _24434_ (.A(_02375_),
    .B(_20244_),
    .Y(_20245_));
 sky130_fd_sc_hd__nand2_1 _24435_ (.A(net350),
    .B(_19796_),
    .Y(_20246_));
 sky130_fd_sc_hd__nand2_1 _24436_ (.A(_20245_),
    .B(_20246_),
    .Y(_20247_));
 sky130_fd_sc_hd__nor2_1 _24437_ (.A(_19431_),
    .B(_19793_),
    .Y(_20248_));
 sky130_fd_sc_hd__inv_2 _24438_ (.A(net353),
    .Y(_02384_));
 sky130_vsdinv _24439_ (.A(net321),
    .Y(_20249_));
 sky130_fd_sc_hd__nor2_1 _24440_ (.A(_02384_),
    .B(_20249_),
    .Y(_20250_));
 sky130_fd_sc_hd__or2_1 _24441_ (.A(_20248_),
    .B(_20250_),
    .X(_20251_));
 sky130_fd_sc_hd__nor2_2 _24442_ (.A(_19433_),
    .B(_19795_),
    .Y(_20252_));
 sky130_fd_sc_hd__inv_2 _24443_ (.A(net351),
    .Y(_02378_));
 sky130_vsdinv _24444_ (.A(_19795_),
    .Y(_20253_));
 sky130_fd_sc_hd__nor2_2 _24445_ (.A(_02378_),
    .B(_20253_),
    .Y(_20254_));
 sky130_fd_sc_hd__nor2_4 _24446_ (.A(_20252_),
    .B(_20254_),
    .Y(_20255_));
 sky130_vsdinv _24447_ (.A(_20255_),
    .Y(_20256_));
 sky130_fd_sc_hd__o2111a_1 _24448_ (.A1(_20241_),
    .A2(_20243_),
    .B1(_20247_),
    .C1(_20251_),
    .D1(_20256_),
    .X(_20257_));
 sky130_fd_sc_hd__nor2_2 _24449_ (.A(_19435_),
    .B(_19799_),
    .Y(_20258_));
 sky130_fd_sc_hd__inv_2 _24450_ (.A(net347),
    .Y(_02369_));
 sky130_vsdinv _24451_ (.A(_19799_),
    .Y(_20259_));
 sky130_fd_sc_hd__nor2_2 _24452_ (.A(_02369_),
    .B(_20259_),
    .Y(_20260_));
 sky130_fd_sc_hd__nor2_2 _24453_ (.A(_19436_),
    .B(_19801_),
    .Y(_20261_));
 sky130_fd_sc_hd__inv_2 _24454_ (.A(_19436_),
    .Y(_02363_));
 sky130_vsdinv _24455_ (.A(net313),
    .Y(_20262_));
 sky130_fd_sc_hd__nor2_1 _24456_ (.A(_02363_),
    .B(_20262_),
    .Y(_20263_));
 sky130_fd_sc_hd__o22a_1 _24457_ (.A1(_20258_),
    .A2(_20260_),
    .B1(_20261_),
    .B2(_20263_),
    .X(_20264_));
 sky130_fd_sc_hd__nor2_1 _24458_ (.A(net346),
    .B(_19800_),
    .Y(_20265_));
 sky130_fd_sc_hd__inv_2 _24459_ (.A(net346),
    .Y(_02366_));
 sky130_vsdinv _24460_ (.A(net314),
    .Y(_20266_));
 sky130_fd_sc_hd__nor2_1 _24461_ (.A(_02366_),
    .B(_20266_),
    .Y(_20267_));
 sky130_fd_sc_hd__nor2_2 _24462_ (.A(_20265_),
    .B(_20267_),
    .Y(_20268_));
 sky130_fd_sc_hd__nor2_1 _24463_ (.A(net348),
    .B(_19797_),
    .Y(_20269_));
 sky130_fd_sc_hd__inv_2 _24464_ (.A(net348),
    .Y(_02372_));
 sky130_vsdinv _24465_ (.A(net316),
    .Y(_20270_));
 sky130_fd_sc_hd__nor2_1 _24466_ (.A(_02372_),
    .B(_20270_),
    .Y(_20271_));
 sky130_fd_sc_hd__nor2_2 _24467_ (.A(_20269_),
    .B(_20271_),
    .Y(_20272_));
 sky130_fd_sc_hd__nor2_1 _24468_ (.A(_20268_),
    .B(_20272_),
    .Y(_20273_));
 sky130_fd_sc_hd__and3_1 _24469_ (.A(_20257_),
    .B(_20264_),
    .C(_20273_),
    .X(_20274_));
 sky130_fd_sc_hd__nand2_2 _24470_ (.A(_20240_),
    .B(_20274_),
    .Y(_20275_));
 sky130_fd_sc_hd__nor2_1 _24471_ (.A(net226),
    .B(_19815_),
    .Y(_20276_));
 sky130_vsdinv _24472_ (.A(net332),
    .Y(_20277_));
 sky130_fd_sc_hd__nor2_1 _24473_ (.A(_20110_),
    .B(_20277_),
    .Y(_20278_));
 sky130_fd_sc_hd__or2_1 _24474_ (.A(_20276_),
    .B(_20278_),
    .X(_20279_));
 sky130_fd_sc_hd__nor2_1 _24475_ (.A(net227),
    .B(_19814_),
    .Y(_20280_));
 sky130_fd_sc_hd__nand2_1 _24476_ (.A(net227),
    .B(_19814_),
    .Y(_20281_));
 sky130_fd_sc_hd__or2b_1 _24477_ (.A(_20280_),
    .B_N(_20281_),
    .X(_20282_));
 sky130_fd_sc_hd__nand2_1 _24478_ (.A(_20279_),
    .B(_20282_),
    .Y(_20283_));
 sky130_fd_sc_hd__nor2_2 _24479_ (.A(net225),
    .B(_19816_),
    .Y(_20284_));
 sky130_vsdinv _24480_ (.A(_19816_),
    .Y(_20285_));
 sky130_fd_sc_hd__nor2_1 _24481_ (.A(_20112_),
    .B(_20285_),
    .Y(_20286_));
 sky130_fd_sc_hd__nor2_1 _24482_ (.A(net222),
    .B(_19817_),
    .Y(_20287_));
 sky130_vsdinv _24483_ (.A(net328),
    .Y(_20288_));
 sky130_fd_sc_hd__nor2_1 _24484_ (.A(_20116_),
    .B(_20288_),
    .Y(_20289_));
 sky130_fd_sc_hd__or2_1 _24485_ (.A(_20287_),
    .B(_20289_),
    .X(_20290_));
 sky130_fd_sc_hd__o21ai_1 _24486_ (.A1(_20284_),
    .A2(_20286_),
    .B1(_20290_),
    .Y(_20291_));
 sky130_fd_sc_hd__or2_1 _24487_ (.A(_20283_),
    .B(_20291_),
    .X(_20292_));
 sky130_fd_sc_hd__nor2_1 _24488_ (.A(net339),
    .B(_19808_),
    .Y(_20293_));
 sky130_fd_sc_hd__inv_2 _24489_ (.A(net339),
    .Y(_02345_));
 sky130_vsdinv _24490_ (.A(net307),
    .Y(_20294_));
 sky130_fd_sc_hd__nor2_1 _24491_ (.A(_02345_),
    .B(_20294_),
    .Y(_20295_));
 sky130_fd_sc_hd__nor2_2 _24492_ (.A(_20293_),
    .B(_20295_),
    .Y(_20296_));
 sky130_fd_sc_hd__nor2_1 _24493_ (.A(_19445_),
    .B(_19810_),
    .Y(_20297_));
 sky130_fd_sc_hd__inv_2 _24494_ (.A(net368),
    .Y(_02339_));
 sky130_vsdinv _24495_ (.A(net336),
    .Y(_20298_));
 sky130_fd_sc_hd__nor2_1 _24496_ (.A(_02339_),
    .B(_20298_),
    .Y(_20299_));
 sky130_fd_sc_hd__nor2_1 _24497_ (.A(_20297_),
    .B(_20299_),
    .Y(_20300_));
 sky130_fd_sc_hd__nor2_1 _24498_ (.A(net340),
    .B(_19807_),
    .Y(_20301_));
 sky130_fd_sc_hd__inv_2 _24499_ (.A(net340),
    .Y(_02348_));
 sky130_vsdinv _24500_ (.A(net308),
    .Y(_20302_));
 sky130_fd_sc_hd__nor2_1 _24501_ (.A(_02348_),
    .B(_20302_),
    .Y(_20303_));
 sky130_fd_sc_hd__nor2_2 _24502_ (.A(_20301_),
    .B(_20303_),
    .Y(_20304_));
 sky130_fd_sc_hd__inv_2 _24503_ (.A(net369),
    .Y(_02342_));
 sky130_vsdinv _24504_ (.A(net337),
    .Y(_20305_));
 sky130_fd_sc_hd__nand2_1 _24505_ (.A(_02342_),
    .B(_20305_),
    .Y(_20306_));
 sky130_fd_sc_hd__nand2_1 _24506_ (.A(_19444_),
    .B(_19809_),
    .Y(_20307_));
 sky130_fd_sc_hd__nand2_1 _24507_ (.A(_20306_),
    .B(_20307_),
    .Y(_20308_));
 sky130_vsdinv _24508_ (.A(_20308_),
    .Y(_20309_));
 sky130_fd_sc_hd__or4_4 _24509_ (.A(_20296_),
    .B(_20300_),
    .C(_20304_),
    .D(_20309_),
    .X(_20310_));
 sky130_fd_sc_hd__nor2_1 _24510_ (.A(_19440_),
    .B(_19804_),
    .Y(_20311_));
 sky130_fd_sc_hd__inv_2 _24511_ (.A(net342),
    .Y(_02354_));
 sky130_vsdinv _24512_ (.A(net310),
    .Y(_20312_));
 sky130_fd_sc_hd__nor2_1 _24513_ (.A(_02354_),
    .B(_20312_),
    .Y(_20313_));
 sky130_fd_sc_hd__nor2_2 _24514_ (.A(_20311_),
    .B(_20313_),
    .Y(_20314_));
 sky130_fd_sc_hd__inv_2 _24515_ (.A(_19438_),
    .Y(_02357_));
 sky130_vsdinv _24516_ (.A(net311),
    .Y(_20315_));
 sky130_fd_sc_hd__nand2_1 _24517_ (.A(_02357_),
    .B(_20315_),
    .Y(_20316_));
 sky130_fd_sc_hd__nand2_1 _24518_ (.A(_19438_),
    .B(_19803_),
    .Y(_20317_));
 sky130_fd_sc_hd__nand2_1 _24519_ (.A(_20316_),
    .B(_20317_),
    .Y(_20318_));
 sky130_vsdinv _24520_ (.A(_20318_),
    .Y(_20319_));
 sky130_fd_sc_hd__nor2_1 _24521_ (.A(_19437_),
    .B(_19802_),
    .Y(_20320_));
 sky130_fd_sc_hd__inv_2 _24522_ (.A(_19437_),
    .Y(_02360_));
 sky130_vsdinv _24523_ (.A(net312),
    .Y(_20321_));
 sky130_fd_sc_hd__nor2_1 _24524_ (.A(_02360_),
    .B(_20321_),
    .Y(_20322_));
 sky130_fd_sc_hd__or2_1 _24525_ (.A(_20320_),
    .B(_20322_),
    .X(_20323_));
 sky130_fd_sc_hd__nor2_1 _24526_ (.A(_19441_),
    .B(_19806_),
    .Y(_20324_));
 sky130_fd_sc_hd__inv_2 _24527_ (.A(net341),
    .Y(_02351_));
 sky130_vsdinv _24528_ (.A(net309),
    .Y(_20325_));
 sky130_fd_sc_hd__nor2_1 _24529_ (.A(_02351_),
    .B(_20325_),
    .Y(_20326_));
 sky130_fd_sc_hd__or2_1 _24530_ (.A(_20324_),
    .B(_20326_),
    .X(_20327_));
 sky130_fd_sc_hd__nand2_1 _24531_ (.A(_20323_),
    .B(_20327_),
    .Y(_20328_));
 sky130_fd_sc_hd__or3_4 _24532_ (.A(_20314_),
    .B(_20319_),
    .C(_20328_),
    .X(_20329_));
 sky130_fd_sc_hd__nor2_1 _24533_ (.A(net228),
    .B(_19813_),
    .Y(_20330_));
 sky130_fd_sc_hd__inv_2 _24534_ (.A(net228),
    .Y(_02333_));
 sky130_vsdinv _24535_ (.A(net334),
    .Y(_20331_));
 sky130_fd_sc_hd__nor2_1 _24536_ (.A(_02333_),
    .B(_20331_),
    .Y(_20332_));
 sky130_fd_sc_hd__nor2_2 _24537_ (.A(_20330_),
    .B(_20332_),
    .Y(_20333_));
 sky130_fd_sc_hd__nor2_1 _24538_ (.A(net229),
    .B(_19811_),
    .Y(_20334_));
 sky130_fd_sc_hd__inv_2 _24539_ (.A(net229),
    .Y(_02336_));
 sky130_vsdinv _24540_ (.A(net335),
    .Y(_20335_));
 sky130_fd_sc_hd__nor2_1 _24541_ (.A(_02336_),
    .B(_20335_),
    .Y(_20336_));
 sky130_fd_sc_hd__nor2_2 _24542_ (.A(_20334_),
    .B(_20336_),
    .Y(_20337_));
 sky130_fd_sc_hd__clkinv_4 _24543_ (.A(_19819_),
    .Y(_20338_));
 sky130_fd_sc_hd__nand2_1 _24544_ (.A(_02318_),
    .B(_20338_),
    .Y(_20339_));
 sky130_fd_sc_hd__nand2_1 _24545_ (.A(_19453_),
    .B(_19819_),
    .Y(_20340_));
 sky130_fd_sc_hd__nand2_1 _24546_ (.A(_20339_),
    .B(_20340_),
    .Y(_20341_));
 sky130_fd_sc_hd__or4b_4 _24547_ (.A(_20333_),
    .B(_20337_),
    .C(_02591_),
    .D_N(_20341_),
    .X(_20342_));
 sky130_fd_sc_hd__or4_4 _24548_ (.A(_20292_),
    .B(_20310_),
    .C(_20329_),
    .D(_20342_),
    .X(_20343_));
 sky130_fd_sc_hd__nor2_4 _24549_ (.A(_20275_),
    .B(_20343_),
    .Y(_00000_));
 sky130_fd_sc_hd__and2_1 _24550_ (.A(_18460_),
    .B(_18465_),
    .X(\pcpi_mul.instr_any_mulh ));
 sky130_fd_sc_hd__or3_2 _24551_ (.A(instr_slt),
    .B(instr_slti),
    .C(instr_blt),
    .X(_00006_));
 sky130_fd_sc_hd__or3_2 _24552_ (.A(instr_sltu),
    .B(instr_sltiu),
    .C(instr_bltu),
    .X(_00007_));
 sky130_fd_sc_hd__nand2_1 _24553_ (.A(_18358_),
    .B(_19981_),
    .Y(_00299_));
 sky130_fd_sc_hd__a2111o_1 _24554_ (.A1(_18501_),
    .A2(_00297_),
    .B1(_18311_),
    .C1(_00319_),
    .D1(_00317_),
    .X(_20344_));
 sky130_fd_sc_hd__a21oi_2 _24555_ (.A1(_18324_),
    .A2(_18553_),
    .B1(_20344_),
    .Y(_20345_));
 sky130_fd_sc_hd__or2_1 _24556_ (.A(instr_lhu),
    .B(instr_lh),
    .X(_20346_));
 sky130_fd_sc_hd__a32o_1 _24557_ (.A1(instr_sh),
    .A2(\cpu_state[5] ),
    .A3(_18739_),
    .B1(_18742_),
    .B2(_20346_),
    .X(_20347_));
 sky130_fd_sc_hd__a2bb2o_1 _24558_ (.A1_N(_20132_),
    .A2_N(_20345_),
    .B1(_18741_),
    .B2(_20347_),
    .X(_00047_));
 sky130_fd_sc_hd__clkbuf_4 _24559_ (.A(_20182_),
    .X(_20348_));
 sky130_fd_sc_hd__and3_1 _24560_ (.A(_20195_),
    .B(_20348_),
    .C(_19782_),
    .X(_00336_));
 sky130_fd_sc_hd__o21ai_1 _24561_ (.A1(_18346_),
    .A2(_18312_),
    .B1(_18361_),
    .Y(_00338_));
 sky130_fd_sc_hd__inv_2 _24562_ (.A(alu_eq),
    .Y(_00340_));
 sky130_vsdinv _24563_ (.A(is_slti_blt_slt),
    .Y(_20349_));
 sky130_vsdinv _24564_ (.A(is_sltiu_bltu_sltu),
    .Y(_20350_));
 sky130_fd_sc_hd__and4_1 _24565_ (.A(_18516_),
    .B(_18727_),
    .C(_20349_),
    .D(_20350_),
    .X(_00341_));
 sky130_fd_sc_hd__a22o_1 _24566_ (.A1(is_slti_blt_slt),
    .A2(alu_lts),
    .B1(is_sltiu_bltu_sltu),
    .B2(alu_ltu),
    .X(_20351_));
 sky130_vsdinv _24567_ (.A(alu_ltu),
    .Y(_20352_));
 sky130_vsdinv _24568_ (.A(alu_lts),
    .Y(_20353_));
 sky130_fd_sc_hd__a22o_1 _24569_ (.A1(_20352_),
    .A2(instr_bgeu),
    .B1(instr_bge),
    .B2(_20353_),
    .X(_20354_));
 sky130_fd_sc_hd__a211oi_2 _24570_ (.A1(instr_bne),
    .A2(_00340_),
    .B1(_20351_),
    .C1(_20354_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand2_1 _24571_ (.A(_20895_),
    .B(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__o22ai_1 _24572_ (.A1(_00346_),
    .A2(_20195_),
    .B1(_00339_),
    .B2(_00297_),
    .Y(_00347_));
 sky130_vsdinv _24573_ (.A(_18525_),
    .Y(_20355_));
 sky130_fd_sc_hd__o21a_1 _24574_ (.A1(_19734_),
    .A2(do_waitirq),
    .B1(_20355_),
    .X(_00349_));
 sky130_fd_sc_hd__and2_1 _24575_ (.A(_02410_),
    .B(_00349_),
    .X(_00351_));
 sky130_fd_sc_hd__o21a_1 _24576_ (.A1(_20195_),
    .A2(_18312_),
    .B1(_18498_),
    .X(_00355_));
 sky130_fd_sc_hd__inv_2 _24577_ (.A(\decoded_imm_uj[4] ),
    .Y(_00367_));
 sky130_vsdinv _24578_ (.A(\cpuregs[0][1] ),
    .Y(_00371_));
 sky130_vsdinv _24579_ (.A(\cpuregs[1][1] ),
    .Y(_00372_));
 sky130_vsdinv _24580_ (.A(\cpuregs[2][1] ),
    .Y(_00373_));
 sky130_vsdinv _24581_ (.A(\cpuregs[3][1] ),
    .Y(_00374_));
 sky130_vsdinv _24582_ (.A(\cpuregs[4][1] ),
    .Y(_00376_));
 sky130_vsdinv _24583_ (.A(\cpuregs[5][1] ),
    .Y(_00377_));
 sky130_vsdinv _24584_ (.A(\cpuregs[6][1] ),
    .Y(_00378_));
 sky130_vsdinv _24585_ (.A(\cpuregs[7][1] ),
    .Y(_00379_));
 sky130_vsdinv _24586_ (.A(\cpuregs[8][1] ),
    .Y(_00381_));
 sky130_vsdinv _24587_ (.A(\cpuregs[9][1] ),
    .Y(_00382_));
 sky130_vsdinv _24588_ (.A(\cpuregs[10][1] ),
    .Y(_00383_));
 sky130_vsdinv _24589_ (.A(\cpuregs[11][1] ),
    .Y(_00384_));
 sky130_vsdinv _24590_ (.A(\cpuregs[12][1] ),
    .Y(_00386_));
 sky130_vsdinv _24591_ (.A(\cpuregs[13][1] ),
    .Y(_00387_));
 sky130_vsdinv _24592_ (.A(\cpuregs[14][1] ),
    .Y(_00388_));
 sky130_vsdinv _24593_ (.A(\cpuregs[15][1] ),
    .Y(_00389_));
 sky130_vsdinv _24594_ (.A(\cpuregs[16][1] ),
    .Y(_00392_));
 sky130_vsdinv _24595_ (.A(\cpuregs[17][1] ),
    .Y(_00393_));
 sky130_vsdinv _24596_ (.A(\cpuregs[18][1] ),
    .Y(_00394_));
 sky130_vsdinv _24597_ (.A(\cpuregs[19][1] ),
    .Y(_00395_));
 sky130_vsdinv _24598_ (.A(\cpuregs[0][2] ),
    .Y(_00398_));
 sky130_vsdinv _24599_ (.A(\cpuregs[1][2] ),
    .Y(_00399_));
 sky130_vsdinv _24600_ (.A(\cpuregs[2][2] ),
    .Y(_00400_));
 sky130_vsdinv _24601_ (.A(\cpuregs[3][2] ),
    .Y(_00401_));
 sky130_vsdinv _24602_ (.A(\cpuregs[4][2] ),
    .Y(_00403_));
 sky130_vsdinv _24603_ (.A(\cpuregs[5][2] ),
    .Y(_00404_));
 sky130_vsdinv _24604_ (.A(\cpuregs[6][2] ),
    .Y(_00405_));
 sky130_vsdinv _24605_ (.A(\cpuregs[7][2] ),
    .Y(_00406_));
 sky130_vsdinv _24606_ (.A(\cpuregs[8][2] ),
    .Y(_00408_));
 sky130_vsdinv _24607_ (.A(\cpuregs[9][2] ),
    .Y(_00409_));
 sky130_vsdinv _24608_ (.A(\cpuregs[10][2] ),
    .Y(_00410_));
 sky130_vsdinv _24609_ (.A(\cpuregs[11][2] ),
    .Y(_00411_));
 sky130_vsdinv _24610_ (.A(\cpuregs[12][2] ),
    .Y(_00413_));
 sky130_vsdinv _24611_ (.A(\cpuregs[13][2] ),
    .Y(_00414_));
 sky130_vsdinv _24612_ (.A(\cpuregs[14][2] ),
    .Y(_00415_));
 sky130_vsdinv _24613_ (.A(\cpuregs[15][2] ),
    .Y(_00416_));
 sky130_vsdinv _24614_ (.A(\cpuregs[16][2] ),
    .Y(_00419_));
 sky130_vsdinv _24615_ (.A(\cpuregs[17][2] ),
    .Y(_00420_));
 sky130_vsdinv _24616_ (.A(\cpuregs[18][2] ),
    .Y(_00421_));
 sky130_vsdinv _24617_ (.A(\cpuregs[19][2] ),
    .Y(_00422_));
 sky130_vsdinv _24618_ (.A(\cpuregs[0][3] ),
    .Y(_00425_));
 sky130_vsdinv _24619_ (.A(\cpuregs[1][3] ),
    .Y(_00426_));
 sky130_vsdinv _24620_ (.A(\cpuregs[2][3] ),
    .Y(_00427_));
 sky130_vsdinv _24621_ (.A(\cpuregs[3][3] ),
    .Y(_00428_));
 sky130_vsdinv _24622_ (.A(\cpuregs[4][3] ),
    .Y(_00430_));
 sky130_vsdinv _24623_ (.A(\cpuregs[5][3] ),
    .Y(_00431_));
 sky130_vsdinv _24624_ (.A(\cpuregs[6][3] ),
    .Y(_00432_));
 sky130_vsdinv _24625_ (.A(\cpuregs[7][3] ),
    .Y(_00433_));
 sky130_vsdinv _24626_ (.A(\cpuregs[8][3] ),
    .Y(_00435_));
 sky130_vsdinv _24627_ (.A(\cpuregs[9][3] ),
    .Y(_00436_));
 sky130_vsdinv _24628_ (.A(\cpuregs[10][3] ),
    .Y(_00437_));
 sky130_vsdinv _24629_ (.A(\cpuregs[11][3] ),
    .Y(_00438_));
 sky130_vsdinv _24630_ (.A(\cpuregs[12][3] ),
    .Y(_00440_));
 sky130_vsdinv _24631_ (.A(\cpuregs[13][3] ),
    .Y(_00441_));
 sky130_vsdinv _24632_ (.A(\cpuregs[14][3] ),
    .Y(_00442_));
 sky130_vsdinv _24633_ (.A(\cpuregs[15][3] ),
    .Y(_00443_));
 sky130_vsdinv _24634_ (.A(\cpuregs[16][3] ),
    .Y(_00446_));
 sky130_vsdinv _24635_ (.A(\cpuregs[17][3] ),
    .Y(_00447_));
 sky130_vsdinv _24636_ (.A(\cpuregs[18][3] ),
    .Y(_00448_));
 sky130_vsdinv _24637_ (.A(\cpuregs[19][3] ),
    .Y(_00449_));
 sky130_vsdinv _24638_ (.A(\cpuregs[0][4] ),
    .Y(_00452_));
 sky130_vsdinv _24639_ (.A(\cpuregs[1][4] ),
    .Y(_00453_));
 sky130_vsdinv _24640_ (.A(\cpuregs[2][4] ),
    .Y(_00454_));
 sky130_vsdinv _24641_ (.A(\cpuregs[3][4] ),
    .Y(_00455_));
 sky130_vsdinv _24642_ (.A(\cpuregs[4][4] ),
    .Y(_00457_));
 sky130_vsdinv _24643_ (.A(\cpuregs[5][4] ),
    .Y(_00458_));
 sky130_vsdinv _24644_ (.A(\cpuregs[6][4] ),
    .Y(_00459_));
 sky130_vsdinv _24645_ (.A(\cpuregs[7][4] ),
    .Y(_00460_));
 sky130_vsdinv _24646_ (.A(\cpuregs[8][4] ),
    .Y(_00462_));
 sky130_vsdinv _24647_ (.A(\cpuregs[9][4] ),
    .Y(_00463_));
 sky130_vsdinv _24648_ (.A(\cpuregs[10][4] ),
    .Y(_00464_));
 sky130_vsdinv _24649_ (.A(\cpuregs[11][4] ),
    .Y(_00465_));
 sky130_vsdinv _24650_ (.A(\cpuregs[12][4] ),
    .Y(_00467_));
 sky130_vsdinv _24651_ (.A(\cpuregs[13][4] ),
    .Y(_00468_));
 sky130_vsdinv _24652_ (.A(\cpuregs[14][4] ),
    .Y(_00469_));
 sky130_vsdinv _24653_ (.A(\cpuregs[15][4] ),
    .Y(_00470_));
 sky130_vsdinv _24654_ (.A(\cpuregs[16][4] ),
    .Y(_00473_));
 sky130_vsdinv _24655_ (.A(\cpuregs[17][4] ),
    .Y(_00474_));
 sky130_vsdinv _24656_ (.A(\cpuregs[18][4] ),
    .Y(_00475_));
 sky130_vsdinv _24657_ (.A(\cpuregs[19][4] ),
    .Y(_00476_));
 sky130_vsdinv _24658_ (.A(\cpuregs[0][5] ),
    .Y(_00479_));
 sky130_vsdinv _24659_ (.A(\cpuregs[1][5] ),
    .Y(_00480_));
 sky130_vsdinv _24660_ (.A(\cpuregs[2][5] ),
    .Y(_00481_));
 sky130_vsdinv _24661_ (.A(\cpuregs[3][5] ),
    .Y(_00482_));
 sky130_vsdinv _24662_ (.A(\cpuregs[4][5] ),
    .Y(_00484_));
 sky130_vsdinv _24663_ (.A(\cpuregs[5][5] ),
    .Y(_00485_));
 sky130_vsdinv _24664_ (.A(\cpuregs[6][5] ),
    .Y(_00486_));
 sky130_vsdinv _24665_ (.A(\cpuregs[7][5] ),
    .Y(_00487_));
 sky130_vsdinv _24666_ (.A(\cpuregs[8][5] ),
    .Y(_00489_));
 sky130_vsdinv _24667_ (.A(\cpuregs[9][5] ),
    .Y(_00490_));
 sky130_vsdinv _24668_ (.A(\cpuregs[10][5] ),
    .Y(_00491_));
 sky130_vsdinv _24669_ (.A(\cpuregs[11][5] ),
    .Y(_00492_));
 sky130_vsdinv _24670_ (.A(\cpuregs[12][5] ),
    .Y(_00494_));
 sky130_vsdinv _24671_ (.A(\cpuregs[13][5] ),
    .Y(_00495_));
 sky130_vsdinv _24672_ (.A(\cpuregs[14][5] ),
    .Y(_00496_));
 sky130_vsdinv _24673_ (.A(\cpuregs[15][5] ),
    .Y(_00497_));
 sky130_vsdinv _24674_ (.A(\cpuregs[16][5] ),
    .Y(_00500_));
 sky130_vsdinv _24675_ (.A(\cpuregs[17][5] ),
    .Y(_00501_));
 sky130_vsdinv _24676_ (.A(\cpuregs[18][5] ),
    .Y(_00502_));
 sky130_vsdinv _24677_ (.A(\cpuregs[19][5] ),
    .Y(_00503_));
 sky130_vsdinv _24678_ (.A(\cpuregs[0][6] ),
    .Y(_00506_));
 sky130_vsdinv _24679_ (.A(\cpuregs[1][6] ),
    .Y(_00507_));
 sky130_vsdinv _24680_ (.A(\cpuregs[2][6] ),
    .Y(_00508_));
 sky130_vsdinv _24681_ (.A(\cpuregs[3][6] ),
    .Y(_00509_));
 sky130_vsdinv _24682_ (.A(\cpuregs[4][6] ),
    .Y(_00511_));
 sky130_vsdinv _24683_ (.A(\cpuregs[5][6] ),
    .Y(_00512_));
 sky130_vsdinv _24684_ (.A(\cpuregs[6][6] ),
    .Y(_00513_));
 sky130_vsdinv _24685_ (.A(\cpuregs[7][6] ),
    .Y(_00514_));
 sky130_vsdinv _24686_ (.A(\cpuregs[8][6] ),
    .Y(_00516_));
 sky130_vsdinv _24687_ (.A(\cpuregs[9][6] ),
    .Y(_00517_));
 sky130_vsdinv _24688_ (.A(\cpuregs[10][6] ),
    .Y(_00518_));
 sky130_vsdinv _24689_ (.A(\cpuregs[11][6] ),
    .Y(_00519_));
 sky130_vsdinv _24690_ (.A(\cpuregs[12][6] ),
    .Y(_00521_));
 sky130_vsdinv _24691_ (.A(\cpuregs[13][6] ),
    .Y(_00522_));
 sky130_vsdinv _24692_ (.A(\cpuregs[14][6] ),
    .Y(_00523_));
 sky130_vsdinv _24693_ (.A(\cpuregs[15][6] ),
    .Y(_00524_));
 sky130_vsdinv _24694_ (.A(\cpuregs[16][6] ),
    .Y(_00527_));
 sky130_vsdinv _24695_ (.A(\cpuregs[17][6] ),
    .Y(_00528_));
 sky130_vsdinv _24696_ (.A(\cpuregs[18][6] ),
    .Y(_00529_));
 sky130_vsdinv _24697_ (.A(\cpuregs[19][6] ),
    .Y(_00530_));
 sky130_vsdinv _24698_ (.A(\cpuregs[0][7] ),
    .Y(_00533_));
 sky130_vsdinv _24699_ (.A(\cpuregs[1][7] ),
    .Y(_00534_));
 sky130_vsdinv _24700_ (.A(\cpuregs[2][7] ),
    .Y(_00535_));
 sky130_vsdinv _24701_ (.A(\cpuregs[3][7] ),
    .Y(_00536_));
 sky130_vsdinv _24702_ (.A(\cpuregs[4][7] ),
    .Y(_00538_));
 sky130_vsdinv _24703_ (.A(\cpuregs[5][7] ),
    .Y(_00539_));
 sky130_vsdinv _24704_ (.A(\cpuregs[6][7] ),
    .Y(_00540_));
 sky130_vsdinv _24705_ (.A(\cpuregs[7][7] ),
    .Y(_00541_));
 sky130_vsdinv _24706_ (.A(\cpuregs[8][7] ),
    .Y(_00543_));
 sky130_vsdinv _24707_ (.A(\cpuregs[9][7] ),
    .Y(_00544_));
 sky130_vsdinv _24708_ (.A(\cpuregs[10][7] ),
    .Y(_00545_));
 sky130_vsdinv _24709_ (.A(\cpuregs[11][7] ),
    .Y(_00546_));
 sky130_vsdinv _24710_ (.A(\cpuregs[12][7] ),
    .Y(_00548_));
 sky130_vsdinv _24711_ (.A(\cpuregs[13][7] ),
    .Y(_00549_));
 sky130_vsdinv _24712_ (.A(\cpuregs[14][7] ),
    .Y(_00550_));
 sky130_vsdinv _24713_ (.A(\cpuregs[15][7] ),
    .Y(_00551_));
 sky130_vsdinv _24714_ (.A(\cpuregs[16][7] ),
    .Y(_00554_));
 sky130_vsdinv _24715_ (.A(\cpuregs[17][7] ),
    .Y(_00555_));
 sky130_vsdinv _24716_ (.A(\cpuregs[18][7] ),
    .Y(_00556_));
 sky130_vsdinv _24717_ (.A(\cpuregs[19][7] ),
    .Y(_00557_));
 sky130_vsdinv _24718_ (.A(\cpuregs[0][8] ),
    .Y(_00560_));
 sky130_vsdinv _24719_ (.A(\cpuregs[1][8] ),
    .Y(_00561_));
 sky130_vsdinv _24720_ (.A(\cpuregs[2][8] ),
    .Y(_00562_));
 sky130_vsdinv _24721_ (.A(\cpuregs[3][8] ),
    .Y(_00563_));
 sky130_vsdinv _24722_ (.A(\cpuregs[4][8] ),
    .Y(_00565_));
 sky130_vsdinv _24723_ (.A(\cpuregs[5][8] ),
    .Y(_00566_));
 sky130_vsdinv _24724_ (.A(\cpuregs[6][8] ),
    .Y(_00567_));
 sky130_vsdinv _24725_ (.A(\cpuregs[7][8] ),
    .Y(_00568_));
 sky130_vsdinv _24726_ (.A(\cpuregs[8][8] ),
    .Y(_00570_));
 sky130_vsdinv _24727_ (.A(\cpuregs[9][8] ),
    .Y(_00571_));
 sky130_vsdinv _24728_ (.A(\cpuregs[10][8] ),
    .Y(_00572_));
 sky130_vsdinv _24729_ (.A(\cpuregs[11][8] ),
    .Y(_00573_));
 sky130_vsdinv _24730_ (.A(\cpuregs[12][8] ),
    .Y(_00575_));
 sky130_vsdinv _24731_ (.A(\cpuregs[13][8] ),
    .Y(_00576_));
 sky130_vsdinv _24732_ (.A(\cpuregs[14][8] ),
    .Y(_00577_));
 sky130_vsdinv _24733_ (.A(\cpuregs[15][8] ),
    .Y(_00578_));
 sky130_vsdinv _24734_ (.A(\cpuregs[16][8] ),
    .Y(_00581_));
 sky130_vsdinv _24735_ (.A(\cpuregs[17][8] ),
    .Y(_00582_));
 sky130_vsdinv _24736_ (.A(\cpuregs[18][8] ),
    .Y(_00583_));
 sky130_vsdinv _24737_ (.A(\cpuregs[19][8] ),
    .Y(_00584_));
 sky130_vsdinv _24738_ (.A(\cpuregs[0][9] ),
    .Y(_00587_));
 sky130_vsdinv _24739_ (.A(\cpuregs[1][9] ),
    .Y(_00588_));
 sky130_vsdinv _24740_ (.A(\cpuregs[2][9] ),
    .Y(_00589_));
 sky130_vsdinv _24741_ (.A(\cpuregs[3][9] ),
    .Y(_00590_));
 sky130_vsdinv _24742_ (.A(\cpuregs[4][9] ),
    .Y(_00592_));
 sky130_vsdinv _24743_ (.A(\cpuregs[5][9] ),
    .Y(_00593_));
 sky130_vsdinv _24744_ (.A(\cpuregs[6][9] ),
    .Y(_00594_));
 sky130_vsdinv _24745_ (.A(\cpuregs[7][9] ),
    .Y(_00595_));
 sky130_vsdinv _24746_ (.A(\cpuregs[8][9] ),
    .Y(_00597_));
 sky130_vsdinv _24747_ (.A(\cpuregs[9][9] ),
    .Y(_00598_));
 sky130_vsdinv _24748_ (.A(\cpuregs[10][9] ),
    .Y(_00599_));
 sky130_vsdinv _24749_ (.A(\cpuregs[11][9] ),
    .Y(_00600_));
 sky130_vsdinv _24750_ (.A(\cpuregs[12][9] ),
    .Y(_00602_));
 sky130_vsdinv _24751_ (.A(\cpuregs[13][9] ),
    .Y(_00603_));
 sky130_vsdinv _24752_ (.A(\cpuregs[14][9] ),
    .Y(_00604_));
 sky130_vsdinv _24753_ (.A(\cpuregs[15][9] ),
    .Y(_00605_));
 sky130_vsdinv _24754_ (.A(\cpuregs[16][9] ),
    .Y(_00608_));
 sky130_vsdinv _24755_ (.A(\cpuregs[17][9] ),
    .Y(_00609_));
 sky130_vsdinv _24756_ (.A(\cpuregs[18][9] ),
    .Y(_00610_));
 sky130_vsdinv _24757_ (.A(\cpuregs[19][9] ),
    .Y(_00611_));
 sky130_vsdinv _24758_ (.A(\cpuregs[0][10] ),
    .Y(_00614_));
 sky130_vsdinv _24759_ (.A(\cpuregs[1][10] ),
    .Y(_00615_));
 sky130_vsdinv _24760_ (.A(\cpuregs[2][10] ),
    .Y(_00616_));
 sky130_vsdinv _24761_ (.A(\cpuregs[3][10] ),
    .Y(_00617_));
 sky130_vsdinv _24762_ (.A(\cpuregs[4][10] ),
    .Y(_00619_));
 sky130_vsdinv _24763_ (.A(\cpuregs[5][10] ),
    .Y(_00620_));
 sky130_vsdinv _24764_ (.A(\cpuregs[6][10] ),
    .Y(_00621_));
 sky130_vsdinv _24765_ (.A(\cpuregs[7][10] ),
    .Y(_00622_));
 sky130_vsdinv _24766_ (.A(\cpuregs[8][10] ),
    .Y(_00624_));
 sky130_vsdinv _24767_ (.A(\cpuregs[9][10] ),
    .Y(_00625_));
 sky130_vsdinv _24768_ (.A(\cpuregs[10][10] ),
    .Y(_00626_));
 sky130_vsdinv _24769_ (.A(\cpuregs[11][10] ),
    .Y(_00627_));
 sky130_vsdinv _24770_ (.A(\cpuregs[12][10] ),
    .Y(_00629_));
 sky130_vsdinv _24771_ (.A(\cpuregs[13][10] ),
    .Y(_00630_));
 sky130_vsdinv _24772_ (.A(\cpuregs[14][10] ),
    .Y(_00631_));
 sky130_vsdinv _24773_ (.A(\cpuregs[15][10] ),
    .Y(_00632_));
 sky130_vsdinv _24774_ (.A(\cpuregs[16][10] ),
    .Y(_00635_));
 sky130_vsdinv _24775_ (.A(\cpuregs[17][10] ),
    .Y(_00636_));
 sky130_vsdinv _24776_ (.A(\cpuregs[18][10] ),
    .Y(_00637_));
 sky130_vsdinv _24777_ (.A(\cpuregs[19][10] ),
    .Y(_00638_));
 sky130_vsdinv _24778_ (.A(\cpuregs[0][11] ),
    .Y(_00641_));
 sky130_vsdinv _24779_ (.A(\cpuregs[1][11] ),
    .Y(_00642_));
 sky130_vsdinv _24780_ (.A(\cpuregs[2][11] ),
    .Y(_00643_));
 sky130_vsdinv _24781_ (.A(\cpuregs[3][11] ),
    .Y(_00644_));
 sky130_vsdinv _24782_ (.A(\cpuregs[4][11] ),
    .Y(_00646_));
 sky130_vsdinv _24783_ (.A(\cpuregs[5][11] ),
    .Y(_00647_));
 sky130_vsdinv _24784_ (.A(\cpuregs[6][11] ),
    .Y(_00648_));
 sky130_vsdinv _24785_ (.A(\cpuregs[7][11] ),
    .Y(_00649_));
 sky130_vsdinv _24786_ (.A(\cpuregs[8][11] ),
    .Y(_00651_));
 sky130_vsdinv _24787_ (.A(\cpuregs[9][11] ),
    .Y(_00652_));
 sky130_vsdinv _24788_ (.A(\cpuregs[10][11] ),
    .Y(_00653_));
 sky130_vsdinv _24789_ (.A(\cpuregs[11][11] ),
    .Y(_00654_));
 sky130_vsdinv _24790_ (.A(\cpuregs[12][11] ),
    .Y(_00656_));
 sky130_vsdinv _24791_ (.A(\cpuregs[13][11] ),
    .Y(_00657_));
 sky130_vsdinv _24792_ (.A(\cpuregs[14][11] ),
    .Y(_00658_));
 sky130_vsdinv _24793_ (.A(\cpuregs[15][11] ),
    .Y(_00659_));
 sky130_vsdinv _24794_ (.A(\cpuregs[16][11] ),
    .Y(_00662_));
 sky130_vsdinv _24795_ (.A(\cpuregs[17][11] ),
    .Y(_00663_));
 sky130_vsdinv _24796_ (.A(\cpuregs[18][11] ),
    .Y(_00664_));
 sky130_vsdinv _24797_ (.A(\cpuregs[19][11] ),
    .Y(_00665_));
 sky130_vsdinv _24798_ (.A(\cpuregs[0][12] ),
    .Y(_00668_));
 sky130_vsdinv _24799_ (.A(\cpuregs[1][12] ),
    .Y(_00669_));
 sky130_vsdinv _24800_ (.A(\cpuregs[2][12] ),
    .Y(_00670_));
 sky130_vsdinv _24801_ (.A(\cpuregs[3][12] ),
    .Y(_00671_));
 sky130_vsdinv _24802_ (.A(\cpuregs[4][12] ),
    .Y(_00673_));
 sky130_vsdinv _24803_ (.A(\cpuregs[5][12] ),
    .Y(_00674_));
 sky130_vsdinv _24804_ (.A(\cpuregs[6][12] ),
    .Y(_00675_));
 sky130_vsdinv _24805_ (.A(\cpuregs[7][12] ),
    .Y(_00676_));
 sky130_vsdinv _24806_ (.A(\cpuregs[8][12] ),
    .Y(_00678_));
 sky130_vsdinv _24807_ (.A(\cpuregs[9][12] ),
    .Y(_00679_));
 sky130_vsdinv _24808_ (.A(\cpuregs[10][12] ),
    .Y(_00680_));
 sky130_vsdinv _24809_ (.A(\cpuregs[11][12] ),
    .Y(_00681_));
 sky130_vsdinv _24810_ (.A(\cpuregs[12][12] ),
    .Y(_00683_));
 sky130_vsdinv _24811_ (.A(\cpuregs[13][12] ),
    .Y(_00684_));
 sky130_vsdinv _24812_ (.A(\cpuregs[14][12] ),
    .Y(_00685_));
 sky130_vsdinv _24813_ (.A(\cpuregs[15][12] ),
    .Y(_00686_));
 sky130_vsdinv _24814_ (.A(\cpuregs[16][12] ),
    .Y(_00689_));
 sky130_vsdinv _24815_ (.A(\cpuregs[17][12] ),
    .Y(_00690_));
 sky130_vsdinv _24816_ (.A(\cpuregs[18][12] ),
    .Y(_00691_));
 sky130_vsdinv _24817_ (.A(\cpuregs[19][12] ),
    .Y(_00692_));
 sky130_vsdinv _24818_ (.A(\cpuregs[0][13] ),
    .Y(_00695_));
 sky130_vsdinv _24819_ (.A(\cpuregs[1][13] ),
    .Y(_00696_));
 sky130_vsdinv _24820_ (.A(\cpuregs[2][13] ),
    .Y(_00697_));
 sky130_vsdinv _24821_ (.A(\cpuregs[3][13] ),
    .Y(_00698_));
 sky130_vsdinv _24822_ (.A(\cpuregs[4][13] ),
    .Y(_00700_));
 sky130_vsdinv _24823_ (.A(\cpuregs[5][13] ),
    .Y(_00701_));
 sky130_vsdinv _24824_ (.A(\cpuregs[6][13] ),
    .Y(_00702_));
 sky130_vsdinv _24825_ (.A(\cpuregs[7][13] ),
    .Y(_00703_));
 sky130_vsdinv _24826_ (.A(\cpuregs[8][13] ),
    .Y(_00705_));
 sky130_vsdinv _24827_ (.A(\cpuregs[9][13] ),
    .Y(_00706_));
 sky130_vsdinv _24828_ (.A(\cpuregs[10][13] ),
    .Y(_00707_));
 sky130_vsdinv _24829_ (.A(\cpuregs[11][13] ),
    .Y(_00708_));
 sky130_vsdinv _24830_ (.A(\cpuregs[12][13] ),
    .Y(_00710_));
 sky130_vsdinv _24831_ (.A(\cpuregs[13][13] ),
    .Y(_00711_));
 sky130_vsdinv _24832_ (.A(\cpuregs[14][13] ),
    .Y(_00712_));
 sky130_vsdinv _24833_ (.A(\cpuregs[15][13] ),
    .Y(_00713_));
 sky130_vsdinv _24834_ (.A(\cpuregs[16][13] ),
    .Y(_00716_));
 sky130_vsdinv _24835_ (.A(\cpuregs[17][13] ),
    .Y(_00717_));
 sky130_vsdinv _24836_ (.A(\cpuregs[18][13] ),
    .Y(_00718_));
 sky130_vsdinv _24837_ (.A(\cpuregs[19][13] ),
    .Y(_00719_));
 sky130_vsdinv _24838_ (.A(\cpuregs[0][14] ),
    .Y(_00722_));
 sky130_vsdinv _24839_ (.A(\cpuregs[1][14] ),
    .Y(_00723_));
 sky130_vsdinv _24840_ (.A(\cpuregs[2][14] ),
    .Y(_00724_));
 sky130_vsdinv _24841_ (.A(\cpuregs[3][14] ),
    .Y(_00725_));
 sky130_vsdinv _24842_ (.A(\cpuregs[4][14] ),
    .Y(_00727_));
 sky130_vsdinv _24843_ (.A(\cpuregs[5][14] ),
    .Y(_00728_));
 sky130_vsdinv _24844_ (.A(\cpuregs[6][14] ),
    .Y(_00729_));
 sky130_vsdinv _24845_ (.A(\cpuregs[7][14] ),
    .Y(_00730_));
 sky130_vsdinv _24846_ (.A(\cpuregs[8][14] ),
    .Y(_00732_));
 sky130_vsdinv _24847_ (.A(\cpuregs[9][14] ),
    .Y(_00733_));
 sky130_vsdinv _24848_ (.A(\cpuregs[10][14] ),
    .Y(_00734_));
 sky130_vsdinv _24849_ (.A(\cpuregs[11][14] ),
    .Y(_00735_));
 sky130_vsdinv _24850_ (.A(\cpuregs[12][14] ),
    .Y(_00737_));
 sky130_vsdinv _24851_ (.A(\cpuregs[13][14] ),
    .Y(_00738_));
 sky130_vsdinv _24852_ (.A(\cpuregs[14][14] ),
    .Y(_00739_));
 sky130_vsdinv _24853_ (.A(\cpuregs[15][14] ),
    .Y(_00740_));
 sky130_vsdinv _24854_ (.A(\cpuregs[16][14] ),
    .Y(_00743_));
 sky130_vsdinv _24855_ (.A(\cpuregs[17][14] ),
    .Y(_00744_));
 sky130_vsdinv _24856_ (.A(\cpuregs[18][14] ),
    .Y(_00745_));
 sky130_vsdinv _24857_ (.A(\cpuregs[19][14] ),
    .Y(_00746_));
 sky130_vsdinv _24858_ (.A(\cpuregs[0][15] ),
    .Y(_00749_));
 sky130_vsdinv _24859_ (.A(\cpuregs[1][15] ),
    .Y(_00750_));
 sky130_vsdinv _24860_ (.A(\cpuregs[2][15] ),
    .Y(_00751_));
 sky130_vsdinv _24861_ (.A(\cpuregs[3][15] ),
    .Y(_00752_));
 sky130_vsdinv _24862_ (.A(\cpuregs[4][15] ),
    .Y(_00754_));
 sky130_vsdinv _24863_ (.A(\cpuregs[5][15] ),
    .Y(_00755_));
 sky130_vsdinv _24864_ (.A(\cpuregs[6][15] ),
    .Y(_00756_));
 sky130_vsdinv _24865_ (.A(\cpuregs[7][15] ),
    .Y(_00757_));
 sky130_vsdinv _24866_ (.A(\cpuregs[8][15] ),
    .Y(_00759_));
 sky130_vsdinv _24867_ (.A(\cpuregs[9][15] ),
    .Y(_00760_));
 sky130_vsdinv _24868_ (.A(\cpuregs[10][15] ),
    .Y(_00761_));
 sky130_vsdinv _24869_ (.A(\cpuregs[11][15] ),
    .Y(_00762_));
 sky130_vsdinv _24870_ (.A(\cpuregs[12][15] ),
    .Y(_00764_));
 sky130_vsdinv _24871_ (.A(\cpuregs[13][15] ),
    .Y(_00765_));
 sky130_vsdinv _24872_ (.A(\cpuregs[14][15] ),
    .Y(_00766_));
 sky130_vsdinv _24873_ (.A(\cpuregs[15][15] ),
    .Y(_00767_));
 sky130_vsdinv _24874_ (.A(\cpuregs[16][15] ),
    .Y(_00770_));
 sky130_vsdinv _24875_ (.A(\cpuregs[17][15] ),
    .Y(_00771_));
 sky130_vsdinv _24876_ (.A(\cpuregs[18][15] ),
    .Y(_00772_));
 sky130_vsdinv _24877_ (.A(\cpuregs[19][15] ),
    .Y(_00773_));
 sky130_vsdinv _24878_ (.A(\cpuregs[0][16] ),
    .Y(_00776_));
 sky130_vsdinv _24879_ (.A(\cpuregs[1][16] ),
    .Y(_00777_));
 sky130_vsdinv _24880_ (.A(\cpuregs[2][16] ),
    .Y(_00778_));
 sky130_vsdinv _24881_ (.A(\cpuregs[3][16] ),
    .Y(_00779_));
 sky130_vsdinv _24882_ (.A(\cpuregs[4][16] ),
    .Y(_00781_));
 sky130_vsdinv _24883_ (.A(\cpuregs[5][16] ),
    .Y(_00782_));
 sky130_vsdinv _24884_ (.A(\cpuregs[6][16] ),
    .Y(_00783_));
 sky130_vsdinv _24885_ (.A(\cpuregs[7][16] ),
    .Y(_00784_));
 sky130_vsdinv _24886_ (.A(\cpuregs[8][16] ),
    .Y(_00786_));
 sky130_vsdinv _24887_ (.A(\cpuregs[9][16] ),
    .Y(_00787_));
 sky130_vsdinv _24888_ (.A(\cpuregs[10][16] ),
    .Y(_00788_));
 sky130_vsdinv _24889_ (.A(\cpuregs[11][16] ),
    .Y(_00789_));
 sky130_vsdinv _24890_ (.A(\cpuregs[12][16] ),
    .Y(_00791_));
 sky130_vsdinv _24891_ (.A(\cpuregs[13][16] ),
    .Y(_00792_));
 sky130_vsdinv _24892_ (.A(\cpuregs[14][16] ),
    .Y(_00793_));
 sky130_vsdinv _24893_ (.A(\cpuregs[15][16] ),
    .Y(_00794_));
 sky130_vsdinv _24894_ (.A(\cpuregs[16][16] ),
    .Y(_00797_));
 sky130_vsdinv _24895_ (.A(\cpuregs[17][16] ),
    .Y(_00798_));
 sky130_vsdinv _24896_ (.A(\cpuregs[18][16] ),
    .Y(_00799_));
 sky130_vsdinv _24897_ (.A(\cpuregs[19][16] ),
    .Y(_00800_));
 sky130_vsdinv _24898_ (.A(\cpuregs[0][17] ),
    .Y(_00803_));
 sky130_vsdinv _24899_ (.A(\cpuregs[1][17] ),
    .Y(_00804_));
 sky130_vsdinv _24900_ (.A(\cpuregs[2][17] ),
    .Y(_00805_));
 sky130_vsdinv _24901_ (.A(\cpuregs[3][17] ),
    .Y(_00806_));
 sky130_vsdinv _24902_ (.A(\cpuregs[4][17] ),
    .Y(_00808_));
 sky130_vsdinv _24903_ (.A(\cpuregs[5][17] ),
    .Y(_00809_));
 sky130_vsdinv _24904_ (.A(\cpuregs[6][17] ),
    .Y(_00810_));
 sky130_vsdinv _24905_ (.A(\cpuregs[7][17] ),
    .Y(_00811_));
 sky130_vsdinv _24906_ (.A(\cpuregs[8][17] ),
    .Y(_00813_));
 sky130_vsdinv _24907_ (.A(\cpuregs[9][17] ),
    .Y(_00814_));
 sky130_vsdinv _24908_ (.A(\cpuregs[10][17] ),
    .Y(_00815_));
 sky130_vsdinv _24909_ (.A(\cpuregs[11][17] ),
    .Y(_00816_));
 sky130_vsdinv _24910_ (.A(\cpuregs[12][17] ),
    .Y(_00818_));
 sky130_vsdinv _24911_ (.A(\cpuregs[13][17] ),
    .Y(_00819_));
 sky130_vsdinv _24912_ (.A(\cpuregs[14][17] ),
    .Y(_00820_));
 sky130_vsdinv _24913_ (.A(\cpuregs[15][17] ),
    .Y(_00821_));
 sky130_vsdinv _24914_ (.A(\cpuregs[16][17] ),
    .Y(_00824_));
 sky130_vsdinv _24915_ (.A(\cpuregs[17][17] ),
    .Y(_00825_));
 sky130_vsdinv _24916_ (.A(\cpuregs[18][17] ),
    .Y(_00826_));
 sky130_vsdinv _24917_ (.A(\cpuregs[19][17] ),
    .Y(_00827_));
 sky130_vsdinv _24918_ (.A(\cpuregs[0][18] ),
    .Y(_00830_));
 sky130_vsdinv _24919_ (.A(\cpuregs[1][18] ),
    .Y(_00831_));
 sky130_vsdinv _24920_ (.A(\cpuregs[2][18] ),
    .Y(_00832_));
 sky130_vsdinv _24921_ (.A(\cpuregs[3][18] ),
    .Y(_00833_));
 sky130_vsdinv _24922_ (.A(\cpuregs[4][18] ),
    .Y(_00835_));
 sky130_vsdinv _24923_ (.A(\cpuregs[5][18] ),
    .Y(_00836_));
 sky130_vsdinv _24924_ (.A(\cpuregs[6][18] ),
    .Y(_00837_));
 sky130_vsdinv _24925_ (.A(\cpuregs[7][18] ),
    .Y(_00838_));
 sky130_vsdinv _24926_ (.A(\cpuregs[8][18] ),
    .Y(_00840_));
 sky130_vsdinv _24927_ (.A(\cpuregs[9][18] ),
    .Y(_00841_));
 sky130_vsdinv _24928_ (.A(\cpuregs[10][18] ),
    .Y(_00842_));
 sky130_vsdinv _24929_ (.A(\cpuregs[11][18] ),
    .Y(_00843_));
 sky130_vsdinv _24930_ (.A(\cpuregs[12][18] ),
    .Y(_00845_));
 sky130_vsdinv _24931_ (.A(\cpuregs[13][18] ),
    .Y(_00846_));
 sky130_vsdinv _24932_ (.A(\cpuregs[14][18] ),
    .Y(_00847_));
 sky130_vsdinv _24933_ (.A(\cpuregs[15][18] ),
    .Y(_00848_));
 sky130_vsdinv _24934_ (.A(\cpuregs[16][18] ),
    .Y(_00851_));
 sky130_vsdinv _24935_ (.A(\cpuregs[17][18] ),
    .Y(_00852_));
 sky130_vsdinv _24936_ (.A(\cpuregs[18][18] ),
    .Y(_00853_));
 sky130_vsdinv _24937_ (.A(\cpuregs[19][18] ),
    .Y(_00854_));
 sky130_vsdinv _24938_ (.A(\cpuregs[0][19] ),
    .Y(_00857_));
 sky130_vsdinv _24939_ (.A(\cpuregs[1][19] ),
    .Y(_00858_));
 sky130_vsdinv _24940_ (.A(\cpuregs[2][19] ),
    .Y(_00859_));
 sky130_vsdinv _24941_ (.A(\cpuregs[3][19] ),
    .Y(_00860_));
 sky130_vsdinv _24942_ (.A(\cpuregs[4][19] ),
    .Y(_00862_));
 sky130_vsdinv _24943_ (.A(\cpuregs[5][19] ),
    .Y(_00863_));
 sky130_vsdinv _24944_ (.A(\cpuregs[6][19] ),
    .Y(_00864_));
 sky130_vsdinv _24945_ (.A(\cpuregs[7][19] ),
    .Y(_00865_));
 sky130_vsdinv _24946_ (.A(\cpuregs[8][19] ),
    .Y(_00867_));
 sky130_vsdinv _24947_ (.A(\cpuregs[9][19] ),
    .Y(_00868_));
 sky130_vsdinv _24948_ (.A(\cpuregs[10][19] ),
    .Y(_00869_));
 sky130_vsdinv _24949_ (.A(\cpuregs[11][19] ),
    .Y(_00870_));
 sky130_vsdinv _24950_ (.A(\cpuregs[12][19] ),
    .Y(_00872_));
 sky130_vsdinv _24951_ (.A(\cpuregs[13][19] ),
    .Y(_00873_));
 sky130_vsdinv _24952_ (.A(\cpuregs[14][19] ),
    .Y(_00874_));
 sky130_vsdinv _24953_ (.A(\cpuregs[15][19] ),
    .Y(_00875_));
 sky130_vsdinv _24954_ (.A(\cpuregs[16][19] ),
    .Y(_00878_));
 sky130_vsdinv _24955_ (.A(\cpuregs[17][19] ),
    .Y(_00879_));
 sky130_vsdinv _24956_ (.A(\cpuregs[18][19] ),
    .Y(_00880_));
 sky130_vsdinv _24957_ (.A(\cpuregs[19][19] ),
    .Y(_00881_));
 sky130_vsdinv _24958_ (.A(\cpuregs[0][20] ),
    .Y(_00884_));
 sky130_vsdinv _24959_ (.A(\cpuregs[1][20] ),
    .Y(_00885_));
 sky130_vsdinv _24960_ (.A(\cpuregs[2][20] ),
    .Y(_00886_));
 sky130_vsdinv _24961_ (.A(\cpuregs[3][20] ),
    .Y(_00887_));
 sky130_vsdinv _24962_ (.A(\cpuregs[4][20] ),
    .Y(_00889_));
 sky130_vsdinv _24963_ (.A(\cpuregs[5][20] ),
    .Y(_00890_));
 sky130_vsdinv _24964_ (.A(\cpuregs[6][20] ),
    .Y(_00891_));
 sky130_vsdinv _24965_ (.A(\cpuregs[7][20] ),
    .Y(_00892_));
 sky130_vsdinv _24966_ (.A(\cpuregs[8][20] ),
    .Y(_00894_));
 sky130_vsdinv _24967_ (.A(\cpuregs[9][20] ),
    .Y(_00895_));
 sky130_vsdinv _24968_ (.A(\cpuregs[10][20] ),
    .Y(_00896_));
 sky130_vsdinv _24969_ (.A(\cpuregs[11][20] ),
    .Y(_00897_));
 sky130_vsdinv _24970_ (.A(\cpuregs[12][20] ),
    .Y(_00899_));
 sky130_vsdinv _24971_ (.A(\cpuregs[13][20] ),
    .Y(_00900_));
 sky130_vsdinv _24972_ (.A(\cpuregs[14][20] ),
    .Y(_00901_));
 sky130_vsdinv _24973_ (.A(\cpuregs[15][20] ),
    .Y(_00902_));
 sky130_vsdinv _24974_ (.A(\cpuregs[16][20] ),
    .Y(_00905_));
 sky130_vsdinv _24975_ (.A(\cpuregs[17][20] ),
    .Y(_00906_));
 sky130_vsdinv _24976_ (.A(\cpuregs[18][20] ),
    .Y(_00907_));
 sky130_vsdinv _24977_ (.A(\cpuregs[19][20] ),
    .Y(_00908_));
 sky130_vsdinv _24978_ (.A(\cpuregs[0][21] ),
    .Y(_00911_));
 sky130_vsdinv _24979_ (.A(\cpuregs[1][21] ),
    .Y(_00912_));
 sky130_vsdinv _24980_ (.A(\cpuregs[2][21] ),
    .Y(_00913_));
 sky130_vsdinv _24981_ (.A(\cpuregs[3][21] ),
    .Y(_00914_));
 sky130_vsdinv _24982_ (.A(\cpuregs[4][21] ),
    .Y(_00916_));
 sky130_vsdinv _24983_ (.A(\cpuregs[5][21] ),
    .Y(_00917_));
 sky130_vsdinv _24984_ (.A(\cpuregs[6][21] ),
    .Y(_00918_));
 sky130_vsdinv _24985_ (.A(\cpuregs[7][21] ),
    .Y(_00919_));
 sky130_vsdinv _24986_ (.A(\cpuregs[8][21] ),
    .Y(_00921_));
 sky130_vsdinv _24987_ (.A(\cpuregs[9][21] ),
    .Y(_00922_));
 sky130_vsdinv _24988_ (.A(\cpuregs[10][21] ),
    .Y(_00923_));
 sky130_vsdinv _24989_ (.A(\cpuregs[11][21] ),
    .Y(_00924_));
 sky130_vsdinv _24990_ (.A(\cpuregs[12][21] ),
    .Y(_00926_));
 sky130_vsdinv _24991_ (.A(\cpuregs[13][21] ),
    .Y(_00927_));
 sky130_vsdinv _24992_ (.A(\cpuregs[14][21] ),
    .Y(_00928_));
 sky130_vsdinv _24993_ (.A(\cpuregs[15][21] ),
    .Y(_00929_));
 sky130_vsdinv _24994_ (.A(\cpuregs[16][21] ),
    .Y(_00932_));
 sky130_vsdinv _24995_ (.A(\cpuregs[17][21] ),
    .Y(_00933_));
 sky130_vsdinv _24996_ (.A(\cpuregs[18][21] ),
    .Y(_00934_));
 sky130_vsdinv _24997_ (.A(\cpuregs[19][21] ),
    .Y(_00935_));
 sky130_vsdinv _24998_ (.A(\cpuregs[0][22] ),
    .Y(_00938_));
 sky130_vsdinv _24999_ (.A(\cpuregs[1][22] ),
    .Y(_00939_));
 sky130_vsdinv _25000_ (.A(\cpuregs[2][22] ),
    .Y(_00940_));
 sky130_vsdinv _25001_ (.A(\cpuregs[3][22] ),
    .Y(_00941_));
 sky130_vsdinv _25002_ (.A(\cpuregs[4][22] ),
    .Y(_00943_));
 sky130_vsdinv _25003_ (.A(\cpuregs[5][22] ),
    .Y(_00944_));
 sky130_vsdinv _25004_ (.A(\cpuregs[6][22] ),
    .Y(_00945_));
 sky130_vsdinv _25005_ (.A(\cpuregs[7][22] ),
    .Y(_00946_));
 sky130_fd_sc_hd__a32o_1 _25006_ (.A1(instr_sw),
    .A2(\cpu_state[5] ),
    .A3(_18739_),
    .B1(_18742_),
    .B2(instr_lw),
    .X(_20356_));
 sky130_fd_sc_hd__nor2_1 _25007_ (.A(_20135_),
    .B(_20345_),
    .Y(_20357_));
 sky130_fd_sc_hd__a211o_1 _25008_ (.A1(_18741_),
    .A2(_20356_),
    .B1(_19370_),
    .C1(_20357_),
    .X(_00045_));
 sky130_vsdinv _25009_ (.A(\cpuregs[8][22] ),
    .Y(_00948_));
 sky130_vsdinv _25010_ (.A(\cpuregs[9][22] ),
    .Y(_00949_));
 sky130_vsdinv _25011_ (.A(\cpuregs[10][22] ),
    .Y(_00950_));
 sky130_vsdinv _25012_ (.A(\cpuregs[11][22] ),
    .Y(_00951_));
 sky130_vsdinv _25013_ (.A(\cpuregs[12][22] ),
    .Y(_00953_));
 sky130_vsdinv _25014_ (.A(\cpuregs[13][22] ),
    .Y(_00954_));
 sky130_vsdinv _25015_ (.A(\cpuregs[14][22] ),
    .Y(_00955_));
 sky130_vsdinv _25016_ (.A(\cpuregs[15][22] ),
    .Y(_00956_));
 sky130_vsdinv _25017_ (.A(\cpuregs[16][22] ),
    .Y(_00959_));
 sky130_vsdinv _25018_ (.A(\cpuregs[17][22] ),
    .Y(_00960_));
 sky130_vsdinv _25019_ (.A(\cpuregs[18][22] ),
    .Y(_00961_));
 sky130_vsdinv _25020_ (.A(\cpuregs[19][22] ),
    .Y(_00962_));
 sky130_vsdinv _25021_ (.A(\cpuregs[0][23] ),
    .Y(_00965_));
 sky130_vsdinv _25022_ (.A(\cpuregs[1][23] ),
    .Y(_00966_));
 sky130_vsdinv _25023_ (.A(\cpuregs[2][23] ),
    .Y(_00967_));
 sky130_vsdinv _25024_ (.A(\cpuregs[3][23] ),
    .Y(_00968_));
 sky130_vsdinv _25025_ (.A(\cpuregs[4][23] ),
    .Y(_00970_));
 sky130_vsdinv _25026_ (.A(\cpuregs[5][23] ),
    .Y(_00971_));
 sky130_vsdinv _25027_ (.A(\cpuregs[6][23] ),
    .Y(_00972_));
 sky130_vsdinv _25028_ (.A(\cpuregs[7][23] ),
    .Y(_00973_));
 sky130_vsdinv _25029_ (.A(\cpuregs[8][23] ),
    .Y(_00975_));
 sky130_vsdinv _25030_ (.A(\cpuregs[9][23] ),
    .Y(_00976_));
 sky130_vsdinv _25031_ (.A(\cpuregs[10][23] ),
    .Y(_00977_));
 sky130_vsdinv _25032_ (.A(\cpuregs[11][23] ),
    .Y(_00978_));
 sky130_vsdinv _25033_ (.A(\cpuregs[12][23] ),
    .Y(_00980_));
 sky130_vsdinv _25034_ (.A(\cpuregs[13][23] ),
    .Y(_00981_));
 sky130_vsdinv _25035_ (.A(\cpuregs[14][23] ),
    .Y(_00982_));
 sky130_vsdinv _25036_ (.A(\cpuregs[15][23] ),
    .Y(_00983_));
 sky130_vsdinv _25037_ (.A(\cpuregs[16][23] ),
    .Y(_00986_));
 sky130_vsdinv _25038_ (.A(\cpuregs[17][23] ),
    .Y(_00987_));
 sky130_vsdinv _25039_ (.A(\cpuregs[18][23] ),
    .Y(_00988_));
 sky130_vsdinv _25040_ (.A(\cpuregs[19][23] ),
    .Y(_00989_));
 sky130_vsdinv _25041_ (.A(\cpuregs[0][24] ),
    .Y(_00992_));
 sky130_vsdinv _25042_ (.A(\cpuregs[1][24] ),
    .Y(_00993_));
 sky130_vsdinv _25043_ (.A(\cpuregs[2][24] ),
    .Y(_00994_));
 sky130_vsdinv _25044_ (.A(\cpuregs[3][24] ),
    .Y(_00995_));
 sky130_vsdinv _25045_ (.A(\cpuregs[4][24] ),
    .Y(_00997_));
 sky130_vsdinv _25046_ (.A(\cpuregs[5][24] ),
    .Y(_00998_));
 sky130_vsdinv _25047_ (.A(\cpuregs[6][24] ),
    .Y(_00999_));
 sky130_vsdinv _25048_ (.A(\cpuregs[7][24] ),
    .Y(_01000_));
 sky130_vsdinv _25049_ (.A(\cpuregs[8][24] ),
    .Y(_01002_));
 sky130_vsdinv _25050_ (.A(\cpuregs[9][24] ),
    .Y(_01003_));
 sky130_vsdinv _25051_ (.A(\cpuregs[10][24] ),
    .Y(_01004_));
 sky130_vsdinv _25052_ (.A(\cpuregs[11][24] ),
    .Y(_01005_));
 sky130_vsdinv _25053_ (.A(\cpuregs[12][24] ),
    .Y(_01007_));
 sky130_vsdinv _25054_ (.A(\cpuregs[13][24] ),
    .Y(_01008_));
 sky130_vsdinv _25055_ (.A(\cpuregs[14][24] ),
    .Y(_01009_));
 sky130_vsdinv _25056_ (.A(\cpuregs[15][24] ),
    .Y(_01010_));
 sky130_vsdinv _25057_ (.A(\cpuregs[16][24] ),
    .Y(_01013_));
 sky130_vsdinv _25058_ (.A(\cpuregs[17][24] ),
    .Y(_01014_));
 sky130_vsdinv _25059_ (.A(\cpuregs[18][24] ),
    .Y(_01015_));
 sky130_vsdinv _25060_ (.A(\cpuregs[19][24] ),
    .Y(_01016_));
 sky130_vsdinv _25061_ (.A(\cpuregs[0][25] ),
    .Y(_01019_));
 sky130_vsdinv _25062_ (.A(\cpuregs[1][25] ),
    .Y(_01020_));
 sky130_vsdinv _25063_ (.A(\cpuregs[2][25] ),
    .Y(_01021_));
 sky130_vsdinv _25064_ (.A(\cpuregs[3][25] ),
    .Y(_01022_));
 sky130_vsdinv _25065_ (.A(\cpuregs[4][25] ),
    .Y(_01024_));
 sky130_vsdinv _25066_ (.A(\cpuregs[5][25] ),
    .Y(_01025_));
 sky130_vsdinv _25067_ (.A(\cpuregs[6][25] ),
    .Y(_01026_));
 sky130_vsdinv _25068_ (.A(\cpuregs[7][25] ),
    .Y(_01027_));
 sky130_fd_sc_hd__nor2_2 _25069_ (.A(\mem_state[1] ),
    .B(_18315_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _25070_ (.A(_18358_),
    .B(_00289_),
    .Y(_00298_));
 sky130_vsdinv _25071_ (.A(\cpuregs[8][25] ),
    .Y(_01029_));
 sky130_vsdinv _25072_ (.A(\cpuregs[9][25] ),
    .Y(_01030_));
 sky130_vsdinv _25073_ (.A(\cpuregs[10][25] ),
    .Y(_01031_));
 sky130_vsdinv _25074_ (.A(\cpuregs[11][25] ),
    .Y(_01032_));
 sky130_vsdinv _25075_ (.A(\cpuregs[12][25] ),
    .Y(_01034_));
 sky130_vsdinv _25076_ (.A(\cpuregs[13][25] ),
    .Y(_01035_));
 sky130_vsdinv _25077_ (.A(\cpuregs[14][25] ),
    .Y(_01036_));
 sky130_vsdinv _25078_ (.A(\cpuregs[15][25] ),
    .Y(_01037_));
 sky130_vsdinv _25079_ (.A(\cpuregs[16][25] ),
    .Y(_01040_));
 sky130_vsdinv _25080_ (.A(\cpuregs[17][25] ),
    .Y(_01041_));
 sky130_vsdinv _25081_ (.A(\cpuregs[18][25] ),
    .Y(_01042_));
 sky130_vsdinv _25082_ (.A(\cpuregs[19][25] ),
    .Y(_01043_));
 sky130_vsdinv _25083_ (.A(\cpuregs[0][26] ),
    .Y(_01046_));
 sky130_vsdinv _25084_ (.A(\cpuregs[1][26] ),
    .Y(_01047_));
 sky130_vsdinv _25085_ (.A(\cpuregs[2][26] ),
    .Y(_01048_));
 sky130_vsdinv _25086_ (.A(\cpuregs[3][26] ),
    .Y(_01049_));
 sky130_vsdinv _25087_ (.A(\cpuregs[4][26] ),
    .Y(_01051_));
 sky130_vsdinv _25088_ (.A(\cpuregs[5][26] ),
    .Y(_01052_));
 sky130_vsdinv _25089_ (.A(\cpuregs[6][26] ),
    .Y(_01053_));
 sky130_vsdinv _25090_ (.A(\cpuregs[7][26] ),
    .Y(_01054_));
 sky130_vsdinv _25091_ (.A(\cpuregs[8][26] ),
    .Y(_01056_));
 sky130_vsdinv _25092_ (.A(\cpuregs[9][26] ),
    .Y(_01057_));
 sky130_vsdinv _25093_ (.A(\cpuregs[10][26] ),
    .Y(_01058_));
 sky130_vsdinv _25094_ (.A(\cpuregs[11][26] ),
    .Y(_01059_));
 sky130_vsdinv _25095_ (.A(\cpuregs[12][26] ),
    .Y(_01061_));
 sky130_vsdinv _25096_ (.A(\cpuregs[13][26] ),
    .Y(_01062_));
 sky130_vsdinv _25097_ (.A(\cpuregs[14][26] ),
    .Y(_01063_));
 sky130_vsdinv _25098_ (.A(\cpuregs[15][26] ),
    .Y(_01064_));
 sky130_vsdinv _25099_ (.A(\cpuregs[16][26] ),
    .Y(_01067_));
 sky130_vsdinv _25100_ (.A(\cpuregs[17][26] ),
    .Y(_01068_));
 sky130_vsdinv _25101_ (.A(\cpuregs[18][26] ),
    .Y(_01069_));
 sky130_vsdinv _25102_ (.A(\cpuregs[19][26] ),
    .Y(_01070_));
 sky130_vsdinv _25103_ (.A(\mem_wordsize[1] ),
    .Y(_20358_));
 sky130_fd_sc_hd__clkbuf_2 _25104_ (.A(_20358_),
    .X(_20359_));
 sky130_fd_sc_hd__clkbuf_2 _25105_ (.A(_18326_),
    .X(_20360_));
 sky130_fd_sc_hd__o211a_1 _25106_ (.A1(instr_lbu),
    .A2(instr_lb),
    .B1(_18334_),
    .C1(_20360_),
    .X(_20361_));
 sky130_fd_sc_hd__a31o_1 _25107_ (.A1(_00291_),
    .A2(instr_sb),
    .A3(\cpu_state[5] ),
    .B1(_20361_),
    .X(_20362_));
 sky130_fd_sc_hd__a2bb2o_1 _25108_ (.A1_N(_20359_),
    .A2_N(_20345_),
    .B1(_18325_),
    .B2(_20362_),
    .X(_00046_));
 sky130_vsdinv _25109_ (.A(\cpuregs[0][27] ),
    .Y(_01073_));
 sky130_vsdinv _25110_ (.A(\cpuregs[1][27] ),
    .Y(_01074_));
 sky130_vsdinv _25111_ (.A(\cpuregs[2][27] ),
    .Y(_01075_));
 sky130_vsdinv _25112_ (.A(\cpuregs[3][27] ),
    .Y(_01076_));
 sky130_vsdinv _25113_ (.A(\cpuregs[4][27] ),
    .Y(_01078_));
 sky130_vsdinv _25114_ (.A(\cpuregs[5][27] ),
    .Y(_01079_));
 sky130_vsdinv _25115_ (.A(\cpuregs[6][27] ),
    .Y(_01080_));
 sky130_vsdinv _25116_ (.A(\cpuregs[7][27] ),
    .Y(_01081_));
 sky130_vsdinv _25117_ (.A(\cpuregs[8][27] ),
    .Y(_01083_));
 sky130_vsdinv _25118_ (.A(\cpuregs[9][27] ),
    .Y(_01084_));
 sky130_vsdinv _25119_ (.A(\cpuregs[10][27] ),
    .Y(_01085_));
 sky130_vsdinv _25120_ (.A(\cpuregs[11][27] ),
    .Y(_01086_));
 sky130_vsdinv _25121_ (.A(\cpuregs[12][27] ),
    .Y(_01088_));
 sky130_vsdinv _25122_ (.A(\cpuregs[13][27] ),
    .Y(_01089_));
 sky130_vsdinv _25123_ (.A(\cpuregs[14][27] ),
    .Y(_01090_));
 sky130_vsdinv _25124_ (.A(\cpuregs[15][27] ),
    .Y(_01091_));
 sky130_vsdinv _25125_ (.A(\cpuregs[16][27] ),
    .Y(_01094_));
 sky130_vsdinv _25126_ (.A(\cpuregs[17][27] ),
    .Y(_01095_));
 sky130_vsdinv _25127_ (.A(\cpuregs[18][27] ),
    .Y(_01096_));
 sky130_vsdinv _25128_ (.A(\cpuregs[19][27] ),
    .Y(_01097_));
 sky130_vsdinv _25129_ (.A(\cpuregs[0][28] ),
    .Y(_01100_));
 sky130_vsdinv _25130_ (.A(\cpuregs[1][28] ),
    .Y(_01101_));
 sky130_vsdinv _25131_ (.A(\cpuregs[2][28] ),
    .Y(_01102_));
 sky130_vsdinv _25132_ (.A(\cpuregs[3][28] ),
    .Y(_01103_));
 sky130_vsdinv _25133_ (.A(\cpuregs[4][28] ),
    .Y(_01105_));
 sky130_vsdinv _25134_ (.A(\cpuregs[5][28] ),
    .Y(_01106_));
 sky130_vsdinv _25135_ (.A(\cpuregs[6][28] ),
    .Y(_01107_));
 sky130_vsdinv _25136_ (.A(\cpuregs[7][28] ),
    .Y(_01108_));
 sky130_vsdinv _25137_ (.A(\cpuregs[8][28] ),
    .Y(_01110_));
 sky130_vsdinv _25138_ (.A(\cpuregs[9][28] ),
    .Y(_01111_));
 sky130_vsdinv _25139_ (.A(\cpuregs[10][28] ),
    .Y(_01112_));
 sky130_vsdinv _25140_ (.A(\cpuregs[11][28] ),
    .Y(_01113_));
 sky130_vsdinv _25141_ (.A(\cpuregs[12][28] ),
    .Y(_01115_));
 sky130_vsdinv _25142_ (.A(\cpuregs[13][28] ),
    .Y(_01116_));
 sky130_vsdinv _25143_ (.A(\cpuregs[14][28] ),
    .Y(_01117_));
 sky130_vsdinv _25144_ (.A(\cpuregs[15][28] ),
    .Y(_01118_));
 sky130_vsdinv _25145_ (.A(\cpuregs[16][28] ),
    .Y(_01121_));
 sky130_vsdinv _25146_ (.A(\cpuregs[17][28] ),
    .Y(_01122_));
 sky130_vsdinv _25147_ (.A(\cpuregs[18][28] ),
    .Y(_01123_));
 sky130_vsdinv _25148_ (.A(\cpuregs[19][28] ),
    .Y(_01124_));
 sky130_vsdinv _25149_ (.A(\cpuregs[0][29] ),
    .Y(_01127_));
 sky130_vsdinv _25150_ (.A(\cpuregs[1][29] ),
    .Y(_01128_));
 sky130_vsdinv _25151_ (.A(\cpuregs[2][29] ),
    .Y(_01129_));
 sky130_vsdinv _25152_ (.A(\cpuregs[3][29] ),
    .Y(_01130_));
 sky130_vsdinv _25153_ (.A(\cpuregs[4][29] ),
    .Y(_01132_));
 sky130_vsdinv _25154_ (.A(\cpuregs[5][29] ),
    .Y(_01133_));
 sky130_vsdinv _25155_ (.A(\cpuregs[6][29] ),
    .Y(_01134_));
 sky130_vsdinv _25156_ (.A(\cpuregs[7][29] ),
    .Y(_01135_));
 sky130_vsdinv _25157_ (.A(\cpuregs[8][29] ),
    .Y(_01137_));
 sky130_vsdinv _25158_ (.A(\cpuregs[9][29] ),
    .Y(_01138_));
 sky130_vsdinv _25159_ (.A(\cpuregs[10][29] ),
    .Y(_01139_));
 sky130_vsdinv _25160_ (.A(\cpuregs[11][29] ),
    .Y(_01140_));
 sky130_vsdinv _25161_ (.A(\cpuregs[12][29] ),
    .Y(_01142_));
 sky130_vsdinv _25162_ (.A(\cpuregs[13][29] ),
    .Y(_01143_));
 sky130_fd_sc_hd__buf_2 _25163_ (.A(latched_branch),
    .X(_20363_));
 sky130_fd_sc_hd__clkbuf_4 _25164_ (.A(_20363_),
    .X(_20364_));
 sky130_fd_sc_hd__and2_1 _25165_ (.A(_20364_),
    .B(_00294_),
    .X(_00295_));
 sky130_vsdinv _25166_ (.A(\cpuregs[14][29] ),
    .Y(_01144_));
 sky130_vsdinv _25167_ (.A(\cpuregs[15][29] ),
    .Y(_01145_));
 sky130_vsdinv _25168_ (.A(\cpuregs[16][29] ),
    .Y(_01148_));
 sky130_vsdinv _25169_ (.A(\cpuregs[17][29] ),
    .Y(_01149_));
 sky130_vsdinv _25170_ (.A(\cpuregs[18][29] ),
    .Y(_01150_));
 sky130_vsdinv _25171_ (.A(\cpuregs[19][29] ),
    .Y(_01151_));
 sky130_vsdinv _25172_ (.A(\cpuregs[0][30] ),
    .Y(_01154_));
 sky130_vsdinv _25173_ (.A(\cpuregs[1][30] ),
    .Y(_01155_));
 sky130_vsdinv _25174_ (.A(\cpuregs[2][30] ),
    .Y(_01156_));
 sky130_vsdinv _25175_ (.A(\cpuregs[3][30] ),
    .Y(_01157_));
 sky130_vsdinv _25176_ (.A(\cpuregs[4][30] ),
    .Y(_01159_));
 sky130_vsdinv _25177_ (.A(\cpuregs[5][30] ),
    .Y(_01160_));
 sky130_vsdinv _25178_ (.A(\cpuregs[6][30] ),
    .Y(_01161_));
 sky130_vsdinv _25179_ (.A(\cpuregs[7][30] ),
    .Y(_01162_));
 sky130_vsdinv _25180_ (.A(\cpuregs[8][30] ),
    .Y(_01164_));
 sky130_vsdinv _25181_ (.A(\cpuregs[9][30] ),
    .Y(_01165_));
 sky130_vsdinv _25182_ (.A(\cpuregs[10][30] ),
    .Y(_01166_));
 sky130_vsdinv _25183_ (.A(\cpuregs[11][30] ),
    .Y(_01167_));
 sky130_vsdinv _25184_ (.A(\cpuregs[12][30] ),
    .Y(_01169_));
 sky130_vsdinv _25185_ (.A(\cpuregs[13][30] ),
    .Y(_01170_));
 sky130_vsdinv _25186_ (.A(\cpuregs[14][30] ),
    .Y(_01171_));
 sky130_vsdinv _25187_ (.A(\cpuregs[15][30] ),
    .Y(_01172_));
 sky130_vsdinv _25188_ (.A(\cpuregs[16][30] ),
    .Y(_01175_));
 sky130_vsdinv _25189_ (.A(\cpuregs[17][30] ),
    .Y(_01176_));
 sky130_vsdinv _25190_ (.A(\cpuregs[18][30] ),
    .Y(_01177_));
 sky130_vsdinv _25191_ (.A(\cpuregs[19][30] ),
    .Y(_01178_));
 sky130_vsdinv _25192_ (.A(\cpuregs[0][31] ),
    .Y(_01181_));
 sky130_vsdinv _25193_ (.A(\cpuregs[1][31] ),
    .Y(_01182_));
 sky130_vsdinv _25194_ (.A(\cpuregs[2][31] ),
    .Y(_01183_));
 sky130_vsdinv _25195_ (.A(\cpuregs[3][31] ),
    .Y(_01184_));
 sky130_vsdinv _25196_ (.A(\cpuregs[4][31] ),
    .Y(_01186_));
 sky130_vsdinv _25197_ (.A(\cpuregs[5][31] ),
    .Y(_01187_));
 sky130_vsdinv _25198_ (.A(\cpuregs[6][31] ),
    .Y(_01188_));
 sky130_vsdinv _25199_ (.A(\cpuregs[7][31] ),
    .Y(_01189_));
 sky130_vsdinv _25200_ (.A(\cpuregs[8][31] ),
    .Y(_01191_));
 sky130_vsdinv _25201_ (.A(\cpuregs[9][31] ),
    .Y(_01192_));
 sky130_vsdinv _25202_ (.A(\cpuregs[10][31] ),
    .Y(_01193_));
 sky130_vsdinv _25203_ (.A(\cpuregs[11][31] ),
    .Y(_01194_));
 sky130_vsdinv _25204_ (.A(\cpuregs[12][31] ),
    .Y(_01196_));
 sky130_vsdinv _25205_ (.A(\cpuregs[13][31] ),
    .Y(_01197_));
 sky130_vsdinv _25206_ (.A(\cpuregs[14][31] ),
    .Y(_01198_));
 sky130_vsdinv _25207_ (.A(\cpuregs[15][31] ),
    .Y(_01199_));
 sky130_vsdinv _25208_ (.A(\cpuregs[16][31] ),
    .Y(_01202_));
 sky130_vsdinv _25209_ (.A(\cpuregs[17][31] ),
    .Y(_01203_));
 sky130_vsdinv _25210_ (.A(\cpuregs[18][31] ),
    .Y(_01204_));
 sky130_vsdinv _25211_ (.A(\cpuregs[19][31] ),
    .Y(_01205_));
 sky130_fd_sc_hd__nor2_1 _25212_ (.A(\timer[5] ),
    .B(\timer[4] ),
    .Y(_20365_));
 sky130_vsdinv _25213_ (.A(_20365_),
    .Y(_20366_));
 sky130_vsdinv _25214_ (.A(\timer[1] ),
    .Y(_20367_));
 sky130_vsdinv _25215_ (.A(\timer[0] ),
    .Y(_20368_));
 sky130_fd_sc_hd__nand2_2 _25216_ (.A(_20367_),
    .B(_20368_),
    .Y(_20369_));
 sky130_fd_sc_hd__or3_4 _25217_ (.A(\timer[3] ),
    .B(\timer[2] ),
    .C(_20369_),
    .X(_20370_));
 sky130_fd_sc_hd__or2_1 _25218_ (.A(_20366_),
    .B(_20370_),
    .X(_20371_));
 sky130_vsdinv _25219_ (.A(_20371_),
    .Y(_20372_));
 sky130_vsdinv _25220_ (.A(\timer[6] ),
    .Y(_20373_));
 sky130_fd_sc_hd__nand2_1 _25221_ (.A(_20372_),
    .B(_20373_),
    .Y(_20374_));
 sky130_fd_sc_hd__nor2_2 _25222_ (.A(\timer[7] ),
    .B(_20374_),
    .Y(_20375_));
 sky130_fd_sc_hd__nor2_1 _25223_ (.A(\timer[9] ),
    .B(\timer[8] ),
    .Y(_20376_));
 sky130_fd_sc_hd__nand2_1 _25224_ (.A(_20375_),
    .B(_20376_),
    .Y(_20377_));
 sky130_fd_sc_hd__nor2_2 _25225_ (.A(\timer[10] ),
    .B(_20377_),
    .Y(_20378_));
 sky130_vsdinv _25226_ (.A(\timer[11] ),
    .Y(_20379_));
 sky130_fd_sc_hd__nor2_1 _25227_ (.A(\timer[13] ),
    .B(\timer[12] ),
    .Y(_20380_));
 sky130_fd_sc_hd__and3_1 _25228_ (.A(_20378_),
    .B(_20379_),
    .C(_20380_),
    .X(_20381_));
 sky130_vsdinv _25229_ (.A(\timer[15] ),
    .Y(_20382_));
 sky130_vsdinv _25230_ (.A(\timer[14] ),
    .Y(_20383_));
 sky130_vsdinv _25231_ (.A(\timer[16] ),
    .Y(_20384_));
 sky130_fd_sc_hd__and3_1 _25232_ (.A(_20382_),
    .B(_20383_),
    .C(_20384_),
    .X(_20385_));
 sky130_fd_sc_hd__nand2_1 _25233_ (.A(_20381_),
    .B(_20385_),
    .Y(_20386_));
 sky130_fd_sc_hd__or2_1 _25234_ (.A(\timer[17] ),
    .B(_20386_),
    .X(_20387_));
 sky130_fd_sc_hd__or2_1 _25235_ (.A(\timer[18] ),
    .B(_20387_),
    .X(_20388_));
 sky130_fd_sc_hd__nor2_1 _25236_ (.A(\timer[19] ),
    .B(_20388_),
    .Y(_20389_));
 sky130_vsdinv _25237_ (.A(\timer[20] ),
    .Y(_20390_));
 sky130_fd_sc_hd__nand2_1 _25238_ (.A(_20389_),
    .B(_20390_),
    .Y(_20391_));
 sky130_fd_sc_hd__or2_1 _25239_ (.A(\timer[21] ),
    .B(_20391_),
    .X(_20392_));
 sky130_fd_sc_hd__or2_1 _25240_ (.A(\timer[22] ),
    .B(_20392_),
    .X(_20393_));
 sky130_fd_sc_hd__nor2_2 _25241_ (.A(\timer[23] ),
    .B(_20393_),
    .Y(_20394_));
 sky130_fd_sc_hd__nor2_1 _25242_ (.A(\timer[25] ),
    .B(\timer[24] ),
    .Y(_20395_));
 sky130_fd_sc_hd__nand2_1 _25243_ (.A(_20394_),
    .B(_20395_),
    .Y(_20396_));
 sky130_fd_sc_hd__or2_2 _25244_ (.A(\timer[26] ),
    .B(_20396_),
    .X(_20397_));
 sky130_fd_sc_hd__nor2_4 _25245_ (.A(\timer[27] ),
    .B(_20397_),
    .Y(_20398_));
 sky130_fd_sc_hd__nor2_1 _25246_ (.A(\timer[29] ),
    .B(\timer[28] ),
    .Y(_20399_));
 sky130_vsdinv _25247_ (.A(\timer[31] ),
    .Y(_20400_));
 sky130_vsdinv _25248_ (.A(\timer[30] ),
    .Y(_20401_));
 sky130_fd_sc_hd__and3_1 _25249_ (.A(_20399_),
    .B(_20400_),
    .C(_20401_),
    .X(_20402_));
 sky130_fd_sc_hd__nand2_4 _25250_ (.A(_20398_),
    .B(_20402_),
    .Y(_20403_));
 sky130_fd_sc_hd__inv_16 _25251_ (.A(_20403_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _25252_ (.A(\timer[0] ),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_1 _25253_ (.A(\timer[1] ),
    .B(\timer[0] ),
    .Y(_20404_));
 sky130_fd_sc_hd__nand2_1 _25254_ (.A(_20369_),
    .B(_20404_),
    .Y(_01211_));
 sky130_vsdinv _25255_ (.A(\timer[2] ),
    .Y(_20405_));
 sky130_fd_sc_hd__xor2_1 _25256_ (.A(_20405_),
    .B(_20369_),
    .X(_01214_));
 sky130_vsdinv _25257_ (.A(\timer[3] ),
    .Y(_20406_));
 sky130_fd_sc_hd__a31o_1 _25258_ (.A1(_20367_),
    .A2(_20368_),
    .A3(_20405_),
    .B1(_20406_),
    .X(_20407_));
 sky130_fd_sc_hd__nand2_1 _25259_ (.A(_20370_),
    .B(_20407_),
    .Y(_01217_));
 sky130_fd_sc_hd__or2_1 _25260_ (.A(\timer[4] ),
    .B(_20370_),
    .X(_20408_));
 sky130_fd_sc_hd__nand2_1 _25261_ (.A(_20370_),
    .B(\timer[4] ),
    .Y(_20409_));
 sky130_fd_sc_hd__nand2_1 _25262_ (.A(_20408_),
    .B(_20409_),
    .Y(_01220_));
 sky130_fd_sc_hd__a21o_1 _25263_ (.A1(_20408_),
    .A2(\timer[5] ),
    .B1(_20372_),
    .X(_01223_));
 sky130_fd_sc_hd__nand2_1 _25264_ (.A(_20371_),
    .B(\timer[6] ),
    .Y(_20410_));
 sky130_fd_sc_hd__nand2_1 _25265_ (.A(_20374_),
    .B(_20410_),
    .Y(_01226_));
 sky130_fd_sc_hd__and2_1 _25266_ (.A(_20374_),
    .B(\timer[7] ),
    .X(_20411_));
 sky130_fd_sc_hd__or2_1 _25267_ (.A(_20375_),
    .B(_20411_),
    .X(_01229_));
 sky130_vsdinv _25268_ (.A(\timer[8] ),
    .Y(_20412_));
 sky130_fd_sc_hd__or2_1 _25269_ (.A(_20412_),
    .B(_20375_),
    .X(_20413_));
 sky130_fd_sc_hd__nand2_1 _25270_ (.A(_20375_),
    .B(_20412_),
    .Y(_20414_));
 sky130_fd_sc_hd__nand2_1 _25271_ (.A(_20413_),
    .B(_20414_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_1 _25272_ (.A(_20414_),
    .B(\timer[9] ),
    .Y(_20415_));
 sky130_fd_sc_hd__nand2_1 _25273_ (.A(_20415_),
    .B(_20377_),
    .Y(_01235_));
 sky130_vsdinv _25274_ (.A(_20378_),
    .Y(_20416_));
 sky130_fd_sc_hd__nand2_1 _25275_ (.A(_20377_),
    .B(\timer[10] ),
    .Y(_20417_));
 sky130_fd_sc_hd__nand2_1 _25276_ (.A(_20416_),
    .B(_20417_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_1 _25277_ (.A(_20416_),
    .B(\timer[11] ),
    .Y(_20418_));
 sky130_fd_sc_hd__nand2_1 _25278_ (.A(_20378_),
    .B(_20379_),
    .Y(_20419_));
 sky130_fd_sc_hd__nand2_1 _25279_ (.A(_20418_),
    .B(_20419_),
    .Y(_01241_));
 sky130_fd_sc_hd__or2_1 _25280_ (.A(\timer[12] ),
    .B(_20419_),
    .X(_20420_));
 sky130_fd_sc_hd__nand2_1 _25281_ (.A(_20419_),
    .B(\timer[12] ),
    .Y(_20421_));
 sky130_fd_sc_hd__nand2_1 _25282_ (.A(_20420_),
    .B(_20421_),
    .Y(_01244_));
 sky130_fd_sc_hd__a21o_1 _25283_ (.A1(_20420_),
    .A2(\timer[13] ),
    .B1(_20381_),
    .X(_01247_));
 sky130_fd_sc_hd__or2_1 _25284_ (.A(_20383_),
    .B(_20381_),
    .X(_20422_));
 sky130_fd_sc_hd__nand2_1 _25285_ (.A(_20381_),
    .B(_20383_),
    .Y(_20423_));
 sky130_fd_sc_hd__nand2_1 _25286_ (.A(_20422_),
    .B(_20423_),
    .Y(_01250_));
 sky130_fd_sc_hd__nor2_1 _25287_ (.A(\timer[15] ),
    .B(_20423_),
    .Y(_20424_));
 sky130_vsdinv _25288_ (.A(_20424_),
    .Y(_20425_));
 sky130_fd_sc_hd__nand2_1 _25289_ (.A(_20423_),
    .B(\timer[15] ),
    .Y(_20426_));
 sky130_fd_sc_hd__nand2_1 _25290_ (.A(_20425_),
    .B(_20426_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_1 _25291_ (.A(_20425_),
    .B(\timer[16] ),
    .Y(_20427_));
 sky130_fd_sc_hd__nand2_1 _25292_ (.A(_20427_),
    .B(_20386_),
    .Y(_01256_));
 sky130_fd_sc_hd__nand2_1 _25293_ (.A(_20386_),
    .B(\timer[17] ),
    .Y(_20428_));
 sky130_fd_sc_hd__nand2_1 _25294_ (.A(_20387_),
    .B(_20428_),
    .Y(_01259_));
 sky130_fd_sc_hd__nand2_1 _25295_ (.A(_20387_),
    .B(\timer[18] ),
    .Y(_20429_));
 sky130_fd_sc_hd__nand2_1 _25296_ (.A(_20388_),
    .B(_20429_),
    .Y(_01262_));
 sky130_fd_sc_hd__and2_1 _25297_ (.A(_20388_),
    .B(\timer[19] ),
    .X(_20430_));
 sky130_fd_sc_hd__or2_1 _25298_ (.A(_20389_),
    .B(_20430_),
    .X(_01265_));
 sky130_fd_sc_hd__or2_1 _25299_ (.A(_20390_),
    .B(_20389_),
    .X(_20431_));
 sky130_fd_sc_hd__nand2_1 _25300_ (.A(_20431_),
    .B(_20391_),
    .Y(_01268_));
 sky130_fd_sc_hd__nand2_1 _25301_ (.A(_20391_),
    .B(\timer[21] ),
    .Y(_20432_));
 sky130_fd_sc_hd__nand2_1 _25302_ (.A(_20392_),
    .B(_20432_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand2_1 _25303_ (.A(_20392_),
    .B(\timer[22] ),
    .Y(_20433_));
 sky130_fd_sc_hd__nand2_1 _25304_ (.A(_20393_),
    .B(_20433_),
    .Y(_01274_));
 sky130_fd_sc_hd__and2_1 _25305_ (.A(_20393_),
    .B(\timer[23] ),
    .X(_20434_));
 sky130_fd_sc_hd__or2_1 _25306_ (.A(_20394_),
    .B(_20434_),
    .X(_01277_));
 sky130_vsdinv _25307_ (.A(\timer[24] ),
    .Y(_20435_));
 sky130_fd_sc_hd__or2_1 _25308_ (.A(_20435_),
    .B(_20394_),
    .X(_20436_));
 sky130_fd_sc_hd__nand2_1 _25309_ (.A(_20394_),
    .B(_20435_),
    .Y(_20437_));
 sky130_fd_sc_hd__nand2_1 _25310_ (.A(_20436_),
    .B(_20437_),
    .Y(_01280_));
 sky130_fd_sc_hd__nand2_1 _25311_ (.A(_20437_),
    .B(\timer[25] ),
    .Y(_20438_));
 sky130_fd_sc_hd__nand2_1 _25312_ (.A(_20438_),
    .B(_20396_),
    .Y(_01283_));
 sky130_fd_sc_hd__nand2_1 _25313_ (.A(_20396_),
    .B(\timer[26] ),
    .Y(_20439_));
 sky130_fd_sc_hd__nand2_1 _25314_ (.A(_20397_),
    .B(_20439_),
    .Y(_01286_));
 sky130_vsdinv _25315_ (.A(_20398_),
    .Y(_20440_));
 sky130_fd_sc_hd__nand2_1 _25316_ (.A(_20397_),
    .B(\timer[27] ),
    .Y(_20441_));
 sky130_fd_sc_hd__nand2_1 _25317_ (.A(_20440_),
    .B(_20441_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_1 _25318_ (.A(_20440_),
    .B(\timer[28] ),
    .Y(_20442_));
 sky130_vsdinv _25319_ (.A(\timer[28] ),
    .Y(_20443_));
 sky130_fd_sc_hd__nand2_1 _25320_ (.A(_20398_),
    .B(_20443_),
    .Y(_20444_));
 sky130_fd_sc_hd__nand2_1 _25321_ (.A(_20442_),
    .B(_20444_),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_1 _25322_ (.A(_20444_),
    .B(\timer[29] ),
    .Y(_20445_));
 sky130_fd_sc_hd__nand2_1 _25323_ (.A(_20398_),
    .B(_20399_),
    .Y(_20446_));
 sky130_fd_sc_hd__nand2_1 _25324_ (.A(_20445_),
    .B(_20446_),
    .Y(_01295_));
 sky130_fd_sc_hd__xor2_1 _25325_ (.A(_20401_),
    .B(_20446_),
    .X(_01298_));
 sky130_fd_sc_hd__a31o_1 _25326_ (.A1(_20398_),
    .A2(_20401_),
    .A3(_20399_),
    .B1(_20400_),
    .X(_20447_));
 sky130_fd_sc_hd__nand2_1 _25327_ (.A(_20447_),
    .B(_20403_),
    .Y(_01301_));
 sky130_fd_sc_hd__buf_4 _25328_ (.A(is_slli_srli_srai),
    .X(_20448_));
 sky130_fd_sc_hd__nor2_8 _25329_ (.A(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .B(_20448_),
    .Y(_01304_));
 sky130_vsdinv _25330_ (.A(\decoded_imm[5] ),
    .Y(_20449_));
 sky130_fd_sc_hd__nor2_1 _25331_ (.A(_20448_),
    .B(_20449_),
    .Y(_01315_));
 sky130_vsdinv _25332_ (.A(\decoded_imm[6] ),
    .Y(_20450_));
 sky130_fd_sc_hd__nor2_1 _25333_ (.A(_20448_),
    .B(_20450_),
    .Y(_01317_));
 sky130_vsdinv _25334_ (.A(\decoded_imm[7] ),
    .Y(_20451_));
 sky130_fd_sc_hd__nor2_1 _25335_ (.A(_20448_),
    .B(_20451_),
    .Y(_01319_));
 sky130_vsdinv _25336_ (.A(\decoded_imm[8] ),
    .Y(_20452_));
 sky130_fd_sc_hd__nor2_1 _25337_ (.A(_20448_),
    .B(_20452_),
    .Y(_01321_));
 sky130_vsdinv _25338_ (.A(\decoded_imm[9] ),
    .Y(_20453_));
 sky130_fd_sc_hd__nor2_1 _25339_ (.A(_20448_),
    .B(_20453_),
    .Y(_01323_));
 sky130_fd_sc_hd__clkbuf_2 _25340_ (.A(_19707_),
    .X(_20454_));
 sky130_vsdinv _25341_ (.A(\decoded_imm[10] ),
    .Y(_20455_));
 sky130_fd_sc_hd__nor2_1 _25342_ (.A(_20454_),
    .B(_20455_),
    .Y(_01325_));
 sky130_vsdinv _25343_ (.A(\decoded_imm[11] ),
    .Y(_20456_));
 sky130_fd_sc_hd__nor2_1 _25344_ (.A(_20454_),
    .B(_20456_),
    .Y(_01327_));
 sky130_vsdinv _25345_ (.A(\decoded_imm[12] ),
    .Y(_20457_));
 sky130_fd_sc_hd__nor2_1 _25346_ (.A(_20454_),
    .B(_20457_),
    .Y(_01329_));
 sky130_vsdinv _25347_ (.A(\decoded_imm[13] ),
    .Y(_20458_));
 sky130_fd_sc_hd__nor2_1 _25348_ (.A(_20454_),
    .B(_20458_),
    .Y(_01331_));
 sky130_vsdinv _25349_ (.A(\decoded_imm[14] ),
    .Y(_20459_));
 sky130_fd_sc_hd__nor2_1 _25350_ (.A(_20454_),
    .B(_20459_),
    .Y(_01333_));
 sky130_vsdinv _25351_ (.A(\decoded_imm[15] ),
    .Y(_20460_));
 sky130_fd_sc_hd__nor2_1 _25352_ (.A(_20454_),
    .B(_20460_),
    .Y(_01335_));
 sky130_fd_sc_hd__clkbuf_2 _25353_ (.A(is_slli_srli_srai),
    .X(_20461_));
 sky130_vsdinv _25354_ (.A(\decoded_imm[16] ),
    .Y(_20462_));
 sky130_fd_sc_hd__nor2_1 _25355_ (.A(_20461_),
    .B(_20462_),
    .Y(_01337_));
 sky130_vsdinv _25356_ (.A(\decoded_imm[17] ),
    .Y(_20463_));
 sky130_fd_sc_hd__nor2_1 _25357_ (.A(_20461_),
    .B(_20463_),
    .Y(_01339_));
 sky130_vsdinv _25358_ (.A(\decoded_imm[18] ),
    .Y(_20464_));
 sky130_fd_sc_hd__nor2_1 _25359_ (.A(_20461_),
    .B(_20464_),
    .Y(_01341_));
 sky130_fd_sc_hd__clkinv_4 _25360_ (.A(\decoded_imm[19] ),
    .Y(_20465_));
 sky130_fd_sc_hd__nor2_1 _25361_ (.A(_20461_),
    .B(_20465_),
    .Y(_01343_));
 sky130_vsdinv _25362_ (.A(\decoded_imm[20] ),
    .Y(_20466_));
 sky130_fd_sc_hd__nor2_1 _25363_ (.A(_20461_),
    .B(_20466_),
    .Y(_01345_));
 sky130_fd_sc_hd__clkinv_4 _25364_ (.A(\decoded_imm[21] ),
    .Y(_20467_));
 sky130_fd_sc_hd__nor2_1 _25365_ (.A(_20461_),
    .B(_20467_),
    .Y(_01347_));
 sky130_fd_sc_hd__clkbuf_2 _25366_ (.A(is_slli_srli_srai),
    .X(_20468_));
 sky130_vsdinv _25367_ (.A(\decoded_imm[22] ),
    .Y(_20469_));
 sky130_fd_sc_hd__nor2_1 _25368_ (.A(_20468_),
    .B(_20469_),
    .Y(_01349_));
 sky130_vsdinv _25369_ (.A(\decoded_imm[23] ),
    .Y(_20470_));
 sky130_fd_sc_hd__nor2_1 _25370_ (.A(_20468_),
    .B(_20470_),
    .Y(_01351_));
 sky130_vsdinv _25371_ (.A(\decoded_imm[24] ),
    .Y(_20471_));
 sky130_fd_sc_hd__nor2_1 _25372_ (.A(_20468_),
    .B(_20471_),
    .Y(_01353_));
 sky130_vsdinv _25373_ (.A(\decoded_imm[25] ),
    .Y(_20472_));
 sky130_fd_sc_hd__nor2_1 _25374_ (.A(_20468_),
    .B(_20472_),
    .Y(_01355_));
 sky130_vsdinv _25375_ (.A(\decoded_imm[26] ),
    .Y(_20473_));
 sky130_fd_sc_hd__nor2_1 _25376_ (.A(_20468_),
    .B(_20473_),
    .Y(_01357_));
 sky130_vsdinv _25377_ (.A(\decoded_imm[27] ),
    .Y(_20474_));
 sky130_fd_sc_hd__nor2_1 _25378_ (.A(_20468_),
    .B(_20474_),
    .Y(_01359_));
 sky130_vsdinv _25379_ (.A(\decoded_imm[28] ),
    .Y(_20475_));
 sky130_fd_sc_hd__nor2_1 _25380_ (.A(_19707_),
    .B(_20475_),
    .Y(_01361_));
 sky130_vsdinv _25381_ (.A(\decoded_imm[29] ),
    .Y(_20476_));
 sky130_fd_sc_hd__nor2_1 _25382_ (.A(_19707_),
    .B(_20476_),
    .Y(_01363_));
 sky130_fd_sc_hd__inv_2 _25383_ (.A(\decoded_imm[30] ),
    .Y(_20477_));
 sky130_fd_sc_hd__nor2_1 _25384_ (.A(_19707_),
    .B(_20477_),
    .Y(_01365_));
 sky130_vsdinv _25385_ (.A(\decoded_imm[31] ),
    .Y(_20478_));
 sky130_fd_sc_hd__nor2_1 _25386_ (.A(_19707_),
    .B(_20478_),
    .Y(_01367_));
 sky130_fd_sc_hd__clkbuf_2 _25387_ (.A(_19776_),
    .X(_20479_));
 sky130_vsdinv _25388_ (.A(\reg_next_pc[0] ),
    .Y(_20480_));
 sky130_fd_sc_hd__nor2_1 _25389_ (.A(_20479_),
    .B(_20480_),
    .Y(_01369_));
 sky130_vsdinv _25390_ (.A(\decoded_imm[0] ),
    .Y(_20481_));
 sky130_fd_sc_hd__nand2_1 _25391_ (.A(_20481_),
    .B(_20119_),
    .Y(_20482_));
 sky130_fd_sc_hd__nand2_1 _25392_ (.A(\decoded_imm[0] ),
    .B(net306),
    .Y(_20483_));
 sky130_fd_sc_hd__and2_1 _25393_ (.A(_20482_),
    .B(_20483_),
    .X(_01371_));
 sky130_fd_sc_hd__nor2_1 _25394_ (.A(_20479_),
    .B(_18867_),
    .Y(_01372_));
 sky130_fd_sc_hd__nor2_1 _25395_ (.A(net317),
    .B(\decoded_imm[1] ),
    .Y(_20484_));
 sky130_fd_sc_hd__nand2_1 _25396_ (.A(_19818_),
    .B(\decoded_imm[1] ),
    .Y(_20485_));
 sky130_fd_sc_hd__or2b_1 _25397_ (.A(_20484_),
    .B_N(_20485_),
    .X(_20486_));
 sky130_fd_sc_hd__xor2_1 _25398_ (.A(_20483_),
    .B(_20486_),
    .X(_01374_));
 sky130_fd_sc_hd__inv_2 _25399_ (.A(\reg_pc[2] ),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_1 _25400_ (.A(_20479_),
    .B(_02073_),
    .Y(_01375_));
 sky130_fd_sc_hd__o21ai_1 _25401_ (.A1(_20483_),
    .A2(_20484_),
    .B1(_20485_),
    .Y(_20487_));
 sky130_fd_sc_hd__xnor2_1 _25402_ (.A(_19817_),
    .B(\decoded_imm[2] ),
    .Y(_20488_));
 sky130_fd_sc_hd__xnor2_1 _25403_ (.A(_20487_),
    .B(_20488_),
    .Y(_01377_));
 sky130_vsdinv _25404_ (.A(\reg_pc[3] ),
    .Y(_20489_));
 sky130_fd_sc_hd__nor2_1 _25405_ (.A(_20479_),
    .B(_20489_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_1 _25406_ (.A(net331),
    .B(\decoded_imm[3] ),
    .Y(_20490_));
 sky130_fd_sc_hd__nand2_1 _25407_ (.A(_19816_),
    .B(\decoded_imm[3] ),
    .Y(_20491_));
 sky130_fd_sc_hd__or2b_1 _25408_ (.A(_20490_),
    .B_N(_20491_),
    .X(_20492_));
 sky130_fd_sc_hd__o21ai_1 _25409_ (.A1(net328),
    .A2(\decoded_imm[2] ),
    .B1(_20487_),
    .Y(_20493_));
 sky130_fd_sc_hd__o21a_1 _25410_ (.A1(_20288_),
    .A2(_20029_),
    .B1(_20493_),
    .X(_20494_));
 sky130_fd_sc_hd__xor2_1 _25411_ (.A(_20492_),
    .B(_20494_),
    .X(_01380_));
 sky130_vsdinv _25412_ (.A(\reg_pc[4] ),
    .Y(_20495_));
 sky130_fd_sc_hd__nor2_1 _25413_ (.A(_20479_),
    .B(_20495_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_1 _25414_ (.A(_19815_),
    .B(\decoded_imm[4] ),
    .Y(_20496_));
 sky130_fd_sc_hd__nor2_2 _25415_ (.A(_20277_),
    .B(_20041_),
    .Y(_20497_));
 sky130_fd_sc_hd__nor2_1 _25416_ (.A(_20496_),
    .B(_20497_),
    .Y(_20498_));
 sky130_fd_sc_hd__o21ai_2 _25417_ (.A1(_20490_),
    .A2(_20494_),
    .B1(_20491_),
    .Y(_20499_));
 sky130_fd_sc_hd__xor2_1 _25418_ (.A(_20498_),
    .B(_20499_),
    .X(_01383_));
 sky130_fd_sc_hd__nor2_1 _25419_ (.A(_20479_),
    .B(_18859_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_1 _25420_ (.A(_19814_),
    .B(\decoded_imm[5] ),
    .Y(_20500_));
 sky130_fd_sc_hd__and2_1 _25421_ (.A(net333),
    .B(\decoded_imm[5] ),
    .X(_20501_));
 sky130_fd_sc_hd__or2_1 _25422_ (.A(_20500_),
    .B(_20501_),
    .X(_20502_));
 sky130_vsdinv _25423_ (.A(_20496_),
    .Y(_20503_));
 sky130_fd_sc_hd__a21oi_4 _25424_ (.A1(_20499_),
    .A2(_20503_),
    .B1(_20497_),
    .Y(_20504_));
 sky130_fd_sc_hd__xor2_1 _25425_ (.A(_20502_),
    .B(_20504_),
    .X(_01386_));
 sky130_fd_sc_hd__clkbuf_2 _25426_ (.A(_19776_),
    .X(_20505_));
 sky130_vsdinv _25427_ (.A(\reg_pc[6] ),
    .Y(_20506_));
 sky130_fd_sc_hd__nor2_1 _25428_ (.A(_20505_),
    .B(_20506_),
    .Y(_01387_));
 sky130_fd_sc_hd__xor2_1 _25429_ (.A(net334),
    .B(\decoded_imm[6] ),
    .X(_20507_));
 sky130_fd_sc_hd__nor2_1 _25430_ (.A(_20500_),
    .B(_20504_),
    .Y(_20508_));
 sky130_fd_sc_hd__or2_1 _25431_ (.A(_20501_),
    .B(_20508_),
    .X(_20509_));
 sky130_fd_sc_hd__or2_1 _25432_ (.A(_20507_),
    .B(_20509_),
    .X(_20510_));
 sky130_fd_sc_hd__nand2_1 _25433_ (.A(_20509_),
    .B(_20507_),
    .Y(_20511_));
 sky130_fd_sc_hd__and2_1 _25434_ (.A(_20510_),
    .B(_20511_),
    .X(_01389_));
 sky130_fd_sc_hd__nor2_1 _25435_ (.A(_20505_),
    .B(_18855_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_1 _25436_ (.A(_19811_),
    .B(\decoded_imm[7] ),
    .Y(_20512_));
 sky130_fd_sc_hd__nor2_1 _25437_ (.A(_20335_),
    .B(_20451_),
    .Y(_20513_));
 sky130_fd_sc_hd__nor2_2 _25438_ (.A(_20512_),
    .B(_20513_),
    .Y(_20514_));
 sky130_fd_sc_hd__o21ai_1 _25439_ (.A1(_20331_),
    .A2(_20450_),
    .B1(_20511_),
    .Y(_20515_));
 sky130_fd_sc_hd__xor2_1 _25440_ (.A(_20514_),
    .B(_20515_),
    .X(_01392_));
 sky130_vsdinv _25441_ (.A(\reg_pc[8] ),
    .Y(_20516_));
 sky130_fd_sc_hd__nor2_1 _25442_ (.A(_20505_),
    .B(_20516_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_1 _25443_ (.A(_19810_),
    .B(\decoded_imm[8] ),
    .Y(_20517_));
 sky130_fd_sc_hd__nor2_1 _25444_ (.A(_20298_),
    .B(_20452_),
    .Y(_20518_));
 sky130_fd_sc_hd__nor2_2 _25445_ (.A(_20517_),
    .B(_20518_),
    .Y(_20519_));
 sky130_fd_sc_hd__and2_1 _25446_ (.A(_20514_),
    .B(_20507_),
    .X(_20520_));
 sky130_fd_sc_hd__o21ai_2 _25447_ (.A1(_20501_),
    .A2(_20508_),
    .B1(_20520_),
    .Y(_20521_));
 sky130_vsdinv _25448_ (.A(_20513_),
    .Y(_20522_));
 sky130_fd_sc_hd__o31a_1 _25449_ (.A1(_20331_),
    .A2(_20450_),
    .A3(_20512_),
    .B1(_20522_),
    .X(_20523_));
 sky130_fd_sc_hd__and2_1 _25450_ (.A(_20521_),
    .B(_20523_),
    .X(_20524_));
 sky130_fd_sc_hd__xnor2_1 _25451_ (.A(_20519_),
    .B(_20524_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor2_1 _25452_ (.A(_20505_),
    .B(_18850_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_1 _25453_ (.A(_19809_),
    .B(\decoded_imm[9] ),
    .Y(_20525_));
 sky130_fd_sc_hd__nor2_1 _25454_ (.A(_20305_),
    .B(_20453_),
    .Y(_20526_));
 sky130_fd_sc_hd__nor2_2 _25455_ (.A(_20525_),
    .B(_20526_),
    .Y(_20527_));
 sky130_vsdinv _25456_ (.A(_20518_),
    .Y(_20528_));
 sky130_fd_sc_hd__o21ai_1 _25457_ (.A1(_20517_),
    .A2(_20524_),
    .B1(_20528_),
    .Y(_20529_));
 sky130_fd_sc_hd__xor2_1 _25458_ (.A(_20527_),
    .B(_20529_),
    .X(_01398_));
 sky130_vsdinv _25459_ (.A(\reg_pc[10] ),
    .Y(_20530_));
 sky130_fd_sc_hd__nor2_1 _25460_ (.A(_20505_),
    .B(_20530_),
    .Y(_01399_));
 sky130_fd_sc_hd__nor2_1 _25461_ (.A(_19808_),
    .B(\decoded_imm[10] ),
    .Y(_20531_));
 sky130_fd_sc_hd__nor2_1 _25462_ (.A(_20294_),
    .B(_20455_),
    .Y(_20532_));
 sky130_fd_sc_hd__or2_1 _25463_ (.A(_20531_),
    .B(_20532_),
    .X(_20533_));
 sky130_vsdinv _25464_ (.A(_20533_),
    .Y(_20534_));
 sky130_fd_sc_hd__o21bai_1 _25465_ (.A1(_20525_),
    .A2(_20528_),
    .B1_N(_20526_),
    .Y(_20535_));
 sky130_fd_sc_hd__nand2_1 _25466_ (.A(_20519_),
    .B(_20527_),
    .Y(_20536_));
 sky130_fd_sc_hd__a21oi_2 _25467_ (.A1(_20521_),
    .A2(_20523_),
    .B1(_20536_),
    .Y(_20537_));
 sky130_fd_sc_hd__or3_2 _25468_ (.A(_20534_),
    .B(_20535_),
    .C(_20537_),
    .X(_20538_));
 sky130_fd_sc_hd__o21bai_2 _25469_ (.A1(_20535_),
    .A2(_20537_),
    .B1_N(_20533_),
    .Y(_20539_));
 sky130_fd_sc_hd__and2_1 _25470_ (.A(_20538_),
    .B(_20539_),
    .X(_01401_));
 sky130_vsdinv _25471_ (.A(\reg_pc[11] ),
    .Y(_20540_));
 sky130_fd_sc_hd__nor2_1 _25472_ (.A(_20505_),
    .B(_20540_),
    .Y(_01402_));
 sky130_vsdinv _25473_ (.A(_20532_),
    .Y(_20541_));
 sky130_fd_sc_hd__nor2_1 _25474_ (.A(_19807_),
    .B(\decoded_imm[11] ),
    .Y(_20542_));
 sky130_fd_sc_hd__nor2_2 _25475_ (.A(_20302_),
    .B(_20456_),
    .Y(_20543_));
 sky130_fd_sc_hd__or2_1 _25476_ (.A(_20542_),
    .B(_20543_),
    .X(_20544_));
 sky130_fd_sc_hd__a21oi_2 _25477_ (.A1(_20539_),
    .A2(_20541_),
    .B1(_20544_),
    .Y(_20545_));
 sky130_fd_sc_hd__and3_1 _25478_ (.A(_20539_),
    .B(_20541_),
    .C(_20544_),
    .X(_20546_));
 sky130_fd_sc_hd__nor2_1 _25479_ (.A(_20545_),
    .B(_20546_),
    .Y(_01404_));
 sky130_fd_sc_hd__clkbuf_2 _25480_ (.A(_19776_),
    .X(_20547_));
 sky130_vsdinv _25481_ (.A(\reg_pc[12] ),
    .Y(_20548_));
 sky130_fd_sc_hd__nor2_1 _25482_ (.A(_20547_),
    .B(_20548_),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_1 _25483_ (.A(net309),
    .B(\decoded_imm[12] ),
    .Y(_20549_));
 sky130_fd_sc_hd__nor2_1 _25484_ (.A(_20325_),
    .B(_20457_),
    .Y(_20550_));
 sky130_fd_sc_hd__or2_1 _25485_ (.A(_20549_),
    .B(_20550_),
    .X(_20551_));
 sky130_vsdinv _25486_ (.A(_20551_),
    .Y(_20552_));
 sky130_fd_sc_hd__or3_2 _25487_ (.A(_20543_),
    .B(_20552_),
    .C(_20545_),
    .X(_20553_));
 sky130_fd_sc_hd__o21bai_2 _25488_ (.A1(_20543_),
    .A2(_20545_),
    .B1_N(_20551_),
    .Y(_20554_));
 sky130_fd_sc_hd__and2_1 _25489_ (.A(_20553_),
    .B(_20554_),
    .X(_01407_));
 sky130_vsdinv _25490_ (.A(\reg_pc[13] ),
    .Y(_20555_));
 sky130_fd_sc_hd__nor2_1 _25491_ (.A(_20547_),
    .B(_20555_),
    .Y(_01408_));
 sky130_vsdinv _25492_ (.A(_20550_),
    .Y(_20556_));
 sky130_fd_sc_hd__nor2_1 _25493_ (.A(_19804_),
    .B(\decoded_imm[13] ),
    .Y(_20557_));
 sky130_fd_sc_hd__nor2_2 _25494_ (.A(_20312_),
    .B(_20458_),
    .Y(_20558_));
 sky130_fd_sc_hd__or2_2 _25495_ (.A(_20557_),
    .B(_20558_),
    .X(_20559_));
 sky130_fd_sc_hd__a21oi_4 _25496_ (.A1(_20554_),
    .A2(_20556_),
    .B1(_20559_),
    .Y(_20560_));
 sky130_fd_sc_hd__and3_1 _25497_ (.A(_20554_),
    .B(_20556_),
    .C(_20559_),
    .X(_20561_));
 sky130_fd_sc_hd__nor2_1 _25498_ (.A(_20560_),
    .B(_20561_),
    .Y(_01410_));
 sky130_vsdinv _25499_ (.A(\reg_pc[14] ),
    .Y(_20562_));
 sky130_fd_sc_hd__nor2_1 _25500_ (.A(_20547_),
    .B(_20562_),
    .Y(_01411_));
 sky130_fd_sc_hd__nor2_1 _25501_ (.A(_19803_),
    .B(\decoded_imm[14] ),
    .Y(_20563_));
 sky130_fd_sc_hd__nor2_1 _25502_ (.A(_20315_),
    .B(_20459_),
    .Y(_20564_));
 sky130_fd_sc_hd__nor2_1 _25503_ (.A(_20563_),
    .B(_20564_),
    .Y(_20565_));
 sky130_fd_sc_hd__or3_2 _25504_ (.A(_20558_),
    .B(_20565_),
    .C(_20560_),
    .X(_20566_));
 sky130_fd_sc_hd__o21ai_2 _25505_ (.A1(_20558_),
    .A2(_20560_),
    .B1(_20565_),
    .Y(_20567_));
 sky130_fd_sc_hd__and2_1 _25506_ (.A(_20566_),
    .B(_20567_),
    .X(_01413_));
 sky130_vsdinv _25507_ (.A(\reg_pc[15] ),
    .Y(_20568_));
 sky130_fd_sc_hd__nor2_1 _25508_ (.A(_20547_),
    .B(_20568_),
    .Y(_01414_));
 sky130_vsdinv _25509_ (.A(_20564_),
    .Y(_20569_));
 sky130_fd_sc_hd__nor2_1 _25510_ (.A(_19802_),
    .B(\decoded_imm[15] ),
    .Y(_20570_));
 sky130_fd_sc_hd__nor2_4 _25511_ (.A(_20321_),
    .B(_20460_),
    .Y(_20571_));
 sky130_fd_sc_hd__nor2_1 _25512_ (.A(_20570_),
    .B(_20571_),
    .Y(_20572_));
 sky130_fd_sc_hd__a21boi_4 _25513_ (.A1(_20567_),
    .A2(_20569_),
    .B1_N(_20572_),
    .Y(_20573_));
 sky130_fd_sc_hd__o211a_1 _25514_ (.A1(_20571_),
    .A2(_20570_),
    .B1(_20569_),
    .C1(_20567_),
    .X(_20574_));
 sky130_fd_sc_hd__nor2_1 _25515_ (.A(_20573_),
    .B(_20574_),
    .Y(_01416_));
 sky130_vsdinv _25516_ (.A(\reg_pc[16] ),
    .Y(_20575_));
 sky130_fd_sc_hd__nor2_1 _25517_ (.A(_20547_),
    .B(_20575_),
    .Y(_01417_));
 sky130_fd_sc_hd__nor2_1 _25518_ (.A(net313),
    .B(\decoded_imm[16] ),
    .Y(_20576_));
 sky130_fd_sc_hd__nor2_1 _25519_ (.A(_20262_),
    .B(_20462_),
    .Y(_20577_));
 sky130_fd_sc_hd__or2_1 _25520_ (.A(_20576_),
    .B(_20577_),
    .X(_20578_));
 sky130_fd_sc_hd__nor2_2 _25521_ (.A(_20571_),
    .B(_20573_),
    .Y(_20579_));
 sky130_fd_sc_hd__xor2_1 _25522_ (.A(_20578_),
    .B(_20579_),
    .X(_01419_));
 sky130_vsdinv _25523_ (.A(\reg_pc[17] ),
    .Y(_20580_));
 sky130_fd_sc_hd__nor2_1 _25524_ (.A(_20547_),
    .B(_20580_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_1 _25525_ (.A(_19800_),
    .B(\decoded_imm[17] ),
    .Y(_20581_));
 sky130_fd_sc_hd__nor2_1 _25526_ (.A(_20266_),
    .B(_20463_),
    .Y(_20582_));
 sky130_fd_sc_hd__nor2_1 _25527_ (.A(_20581_),
    .B(_20582_),
    .Y(_20583_));
 sky130_fd_sc_hd__o21ba_1 _25528_ (.A1(_20576_),
    .A2(_20579_),
    .B1_N(_20577_),
    .X(_20584_));
 sky130_fd_sc_hd__xnor2_1 _25529_ (.A(_20583_),
    .B(_20584_),
    .Y(_01422_));
 sky130_fd_sc_hd__clkbuf_2 _25530_ (.A(instr_lui),
    .X(_20585_));
 sky130_vsdinv _25531_ (.A(\reg_pc[18] ),
    .Y(_20586_));
 sky130_fd_sc_hd__nor2_1 _25532_ (.A(_20585_),
    .B(_20586_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_2 _25533_ (.A(_19799_),
    .B(\decoded_imm[18] ),
    .Y(_20587_));
 sky130_fd_sc_hd__nor2_4 _25534_ (.A(_20259_),
    .B(_20464_),
    .Y(_20588_));
 sky130_fd_sc_hd__nor2_1 _25535_ (.A(_20587_),
    .B(_20588_),
    .Y(_20589_));
 sky130_fd_sc_hd__and2b_1 _25536_ (.A_N(_20578_),
    .B(_20583_),
    .X(_20590_));
 sky130_fd_sc_hd__o21ai_2 _25537_ (.A1(_20571_),
    .A2(_20573_),
    .B1(_20590_),
    .Y(_20591_));
 sky130_vsdinv _25538_ (.A(_20582_),
    .Y(_20592_));
 sky130_fd_sc_hd__o31a_1 _25539_ (.A1(_20262_),
    .A2(_20462_),
    .A3(_20581_),
    .B1(_20592_),
    .X(_20593_));
 sky130_fd_sc_hd__nand2_1 _25540_ (.A(_20591_),
    .B(_20593_),
    .Y(_20594_));
 sky130_fd_sc_hd__xor2_1 _25541_ (.A(_20589_),
    .B(_20594_),
    .X(_01425_));
 sky130_fd_sc_hd__clkinv_4 _25542_ (.A(\reg_pc[19] ),
    .Y(_20595_));
 sky130_fd_sc_hd__nor2_1 _25543_ (.A(_20585_),
    .B(_20595_),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_2 _25544_ (.A(_19797_),
    .B(_20465_),
    .Y(_20596_));
 sky130_fd_sc_hd__nor2_2 _25545_ (.A(\decoded_imm[19] ),
    .B(_20270_),
    .Y(_20597_));
 sky130_fd_sc_hd__a21oi_4 _25546_ (.A1(_20591_),
    .A2(_20593_),
    .B1(_20587_),
    .Y(_20598_));
 sky130_fd_sc_hd__or4_1 _25547_ (.A(_20588_),
    .B(_20596_),
    .C(_20597_),
    .D(_20598_),
    .X(_20599_));
 sky130_fd_sc_hd__o22ai_4 _25548_ (.A1(_20596_),
    .A2(_20597_),
    .B1(_20588_),
    .B2(_20598_),
    .Y(_20600_));
 sky130_fd_sc_hd__and2_1 _25549_ (.A(_20599_),
    .B(_20600_),
    .X(_01428_));
 sky130_vsdinv _25550_ (.A(\reg_pc[20] ),
    .Y(_20601_));
 sky130_fd_sc_hd__nor2_1 _25551_ (.A(_20585_),
    .B(_20601_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_1 _25552_ (.A(_20270_),
    .B(_20465_),
    .Y(_20602_));
 sky130_vsdinv _25553_ (.A(_20602_),
    .Y(_20603_));
 sky130_fd_sc_hd__nor2_1 _25554_ (.A(_19796_),
    .B(\decoded_imm[20] ),
    .Y(_20604_));
 sky130_fd_sc_hd__nor2_4 _25555_ (.A(_20244_),
    .B(_20466_),
    .Y(_20605_));
 sky130_fd_sc_hd__or2_2 _25556_ (.A(_20604_),
    .B(_20605_),
    .X(_20606_));
 sky130_fd_sc_hd__a21oi_4 _25557_ (.A1(_20600_),
    .A2(_20603_),
    .B1(_20606_),
    .Y(_20607_));
 sky130_fd_sc_hd__and3_1 _25558_ (.A(_20600_),
    .B(_20603_),
    .C(_20606_),
    .X(_20608_));
 sky130_fd_sc_hd__nor2_1 _25559_ (.A(_20607_),
    .B(_20608_),
    .Y(_01431_));
 sky130_vsdinv _25560_ (.A(\reg_pc[21] ),
    .Y(_20609_));
 sky130_fd_sc_hd__nor2_1 _25561_ (.A(_20585_),
    .B(_20609_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_2 _25562_ (.A(_19795_),
    .B(_20467_),
    .Y(_20610_));
 sky130_fd_sc_hd__nor2_2 _25563_ (.A(\decoded_imm[21] ),
    .B(_20253_),
    .Y(_20611_));
 sky130_fd_sc_hd__or4_1 _25564_ (.A(_20605_),
    .B(_20610_),
    .C(_20611_),
    .D(_20607_),
    .X(_20612_));
 sky130_fd_sc_hd__o22ai_4 _25565_ (.A1(_20610_),
    .A2(_20611_),
    .B1(_20605_),
    .B2(_20607_),
    .Y(_20613_));
 sky130_fd_sc_hd__and2_1 _25566_ (.A(_20612_),
    .B(_20613_),
    .X(_01434_));
 sky130_vsdinv _25567_ (.A(\reg_pc[22] ),
    .Y(_20614_));
 sky130_fd_sc_hd__nor2_1 _25568_ (.A(_20585_),
    .B(_20614_),
    .Y(_01435_));
 sky130_fd_sc_hd__nor2_1 _25569_ (.A(_20253_),
    .B(_20467_),
    .Y(_20615_));
 sky130_vsdinv _25570_ (.A(_20615_),
    .Y(_20616_));
 sky130_fd_sc_hd__nor2_1 _25571_ (.A(net320),
    .B(\decoded_imm[22] ),
    .Y(_20617_));
 sky130_fd_sc_hd__nor2_4 _25572_ (.A(_20242_),
    .B(_20469_),
    .Y(_20618_));
 sky130_fd_sc_hd__or2_2 _25573_ (.A(_20617_),
    .B(_20618_),
    .X(_20619_));
 sky130_fd_sc_hd__a21oi_4 _25574_ (.A1(_20613_),
    .A2(_20616_),
    .B1(_20619_),
    .Y(_20620_));
 sky130_fd_sc_hd__and3_1 _25575_ (.A(_20613_),
    .B(_20616_),
    .C(_20619_),
    .X(_20621_));
 sky130_fd_sc_hd__nor2_1 _25576_ (.A(_20620_),
    .B(_20621_),
    .Y(_01437_));
 sky130_vsdinv _25577_ (.A(\reg_pc[23] ),
    .Y(_20622_));
 sky130_fd_sc_hd__nor2_1 _25578_ (.A(_20585_),
    .B(_20622_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_2 _25579_ (.A(_19793_),
    .B(_20470_),
    .Y(_20623_));
 sky130_fd_sc_hd__nor2_2 _25580_ (.A(\decoded_imm[23] ),
    .B(_20249_),
    .Y(_20624_));
 sky130_fd_sc_hd__or4_1 _25581_ (.A(_20618_),
    .B(_20623_),
    .C(_20624_),
    .D(_20620_),
    .X(_20625_));
 sky130_fd_sc_hd__o22ai_4 _25582_ (.A1(_20623_),
    .A2(_20624_),
    .B1(_20618_),
    .B2(_20620_),
    .Y(_20626_));
 sky130_fd_sc_hd__and2_1 _25583_ (.A(_20625_),
    .B(_20626_),
    .X(_01440_));
 sky130_fd_sc_hd__clkbuf_2 _25584_ (.A(instr_lui),
    .X(_20627_));
 sky130_vsdinv _25585_ (.A(\reg_pc[24] ),
    .Y(_20628_));
 sky130_fd_sc_hd__nor2_1 _25586_ (.A(_20627_),
    .B(_20628_),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_1 _25587_ (.A(_20217_),
    .B(_20471_),
    .Y(_20629_));
 sky130_fd_sc_hd__nand2_1 _25588_ (.A(_19792_),
    .B(\decoded_imm[24] ),
    .Y(_20630_));
 sky130_fd_sc_hd__nand2_1 _25589_ (.A(_20629_),
    .B(_20630_),
    .Y(_20631_));
 sky130_vsdinv _25590_ (.A(_20631_),
    .Y(_20632_));
 sky130_fd_sc_hd__nand2_1 _25591_ (.A(_19793_),
    .B(\decoded_imm[23] ),
    .Y(_20633_));
 sky130_fd_sc_hd__nand2_1 _25592_ (.A(_20626_),
    .B(_20633_),
    .Y(_20634_));
 sky130_fd_sc_hd__or2_1 _25593_ (.A(_20632_),
    .B(_20634_),
    .X(_20635_));
 sky130_fd_sc_hd__nand2_1 _25594_ (.A(_20634_),
    .B(_20632_),
    .Y(_20636_));
 sky130_fd_sc_hd__and2_1 _25595_ (.A(_20635_),
    .B(_20636_),
    .X(_01443_));
 sky130_vsdinv _25596_ (.A(\reg_pc[25] ),
    .Y(_20637_));
 sky130_fd_sc_hd__nor2_1 _25597_ (.A(_20627_),
    .B(_20637_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _25598_ (.A(_19790_),
    .B(\decoded_imm[25] ),
    .Y(_20638_));
 sky130_fd_sc_hd__nor2_1 _25599_ (.A(_20205_),
    .B(_20472_),
    .Y(_20639_));
 sky130_fd_sc_hd__or2_1 _25600_ (.A(_20638_),
    .B(_20639_),
    .X(_20640_));
 sky130_vsdinv _25601_ (.A(_20640_),
    .Y(_20641_));
 sky130_fd_sc_hd__nand2_1 _25602_ (.A(_20636_),
    .B(_20630_),
    .Y(_20642_));
 sky130_fd_sc_hd__xor2_1 _25603_ (.A(_20641_),
    .B(_20642_),
    .X(_01446_));
 sky130_vsdinv _25604_ (.A(\reg_pc[26] ),
    .Y(_20643_));
 sky130_fd_sc_hd__nor2_1 _25605_ (.A(_20627_),
    .B(_20643_),
    .Y(_01447_));
 sky130_fd_sc_hd__nor2_1 _25606_ (.A(net324),
    .B(\decoded_imm[26] ),
    .Y(_20644_));
 sky130_fd_sc_hd__nor2_4 _25607_ (.A(_20210_),
    .B(_20473_),
    .Y(_20645_));
 sky130_fd_sc_hd__nor2_1 _25608_ (.A(_20644_),
    .B(_20645_),
    .Y(_20646_));
 sky130_fd_sc_hd__o21bai_1 _25609_ (.A1(_20630_),
    .A2(_20638_),
    .B1_N(_20639_),
    .Y(_20647_));
 sky130_fd_sc_hd__nand2_1 _25610_ (.A(_20641_),
    .B(_20632_),
    .Y(_20648_));
 sky130_fd_sc_hd__a21oi_2 _25611_ (.A1(_20626_),
    .A2(_20633_),
    .B1(_20648_),
    .Y(_20649_));
 sky130_fd_sc_hd__or2_1 _25612_ (.A(_20647_),
    .B(_20649_),
    .X(_20650_));
 sky130_fd_sc_hd__nor2_1 _25613_ (.A(_20646_),
    .B(_20650_),
    .Y(_20651_));
 sky130_fd_sc_hd__and2_1 _25614_ (.A(_20650_),
    .B(_20646_),
    .X(_20652_));
 sky130_fd_sc_hd__nor2_1 _25615_ (.A(_20651_),
    .B(_20652_),
    .Y(_01449_));
 sky130_vsdinv _25616_ (.A(\reg_pc[27] ),
    .Y(_20653_));
 sky130_fd_sc_hd__nor2_1 _25617_ (.A(_20627_),
    .B(_20653_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_1 _25618_ (.A(_19789_),
    .B(\decoded_imm[27] ),
    .Y(_20654_));
 sky130_vsdinv _25619_ (.A(_19789_),
    .Y(_20655_));
 sky130_fd_sc_hd__nor2_4 _25620_ (.A(_20655_),
    .B(_20474_),
    .Y(_20656_));
 sky130_fd_sc_hd__nor2_2 _25621_ (.A(_20654_),
    .B(_20656_),
    .Y(_20657_));
 sky130_fd_sc_hd__nor2_1 _25622_ (.A(_20645_),
    .B(_20652_),
    .Y(_20658_));
 sky130_fd_sc_hd__xnor2_1 _25623_ (.A(_20657_),
    .B(_20658_),
    .Y(_01452_));
 sky130_vsdinv _25624_ (.A(\reg_pc[28] ),
    .Y(_20659_));
 sky130_fd_sc_hd__nor2_1 _25625_ (.A(_20627_),
    .B(_20659_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_1 _25626_ (.A(_20646_),
    .B(_20657_),
    .Y(_20660_));
 sky130_fd_sc_hd__o21bai_2 _25627_ (.A1(_20647_),
    .A2(_20649_),
    .B1_N(_20660_),
    .Y(_20661_));
 sky130_vsdinv _25628_ (.A(_20654_),
    .Y(_20662_));
 sky130_fd_sc_hd__a21oi_4 _25629_ (.A1(_20645_),
    .A2(_20662_),
    .B1(_20656_),
    .Y(_20663_));
 sky130_fd_sc_hd__nor2_2 _25630_ (.A(net326),
    .B(\decoded_imm[28] ),
    .Y(_20664_));
 sky130_fd_sc_hd__nor2_4 _25631_ (.A(_20236_),
    .B(_20475_),
    .Y(_20665_));
 sky130_fd_sc_hd__or2_1 _25632_ (.A(_20664_),
    .B(_20665_),
    .X(_20666_));
 sky130_fd_sc_hd__a21oi_1 _25633_ (.A1(_20661_),
    .A2(_20663_),
    .B1(_20666_),
    .Y(_20667_));
 sky130_fd_sc_hd__and3_1 _25634_ (.A(_20661_),
    .B(_20663_),
    .C(_20666_),
    .X(_20668_));
 sky130_fd_sc_hd__nor2_1 _25635_ (.A(_20667_),
    .B(_20668_),
    .Y(_01455_));
 sky130_vsdinv _25636_ (.A(\reg_pc[29] ),
    .Y(_20669_));
 sky130_fd_sc_hd__nor2_1 _25637_ (.A(_20627_),
    .B(_20669_),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_1 _25638_ (.A(_20231_),
    .B(_20476_),
    .Y(_20670_));
 sky130_fd_sc_hd__nand2_2 _25639_ (.A(_19788_),
    .B(\decoded_imm[29] ),
    .Y(_20671_));
 sky130_fd_sc_hd__nand2_1 _25640_ (.A(_20670_),
    .B(_20671_),
    .Y(_20672_));
 sky130_fd_sc_hd__a21oi_4 _25641_ (.A1(_20661_),
    .A2(_20663_),
    .B1(_20664_),
    .Y(_20673_));
 sky130_fd_sc_hd__or3_2 _25642_ (.A(_20665_),
    .B(_20672_),
    .C(_20673_),
    .X(_20674_));
 sky130_fd_sc_hd__o21ai_1 _25643_ (.A1(_20665_),
    .A2(_20673_),
    .B1(_20672_),
    .Y(_20675_));
 sky130_fd_sc_hd__nand2_1 _25644_ (.A(_20674_),
    .B(_20675_),
    .Y(_01458_));
 sky130_vsdinv _25645_ (.A(\reg_pc[30] ),
    .Y(_20676_));
 sky130_fd_sc_hd__nor2_1 _25646_ (.A(_19776_),
    .B(_20676_),
    .Y(_01459_));
 sky130_fd_sc_hd__nor2_1 _25647_ (.A(_19787_),
    .B(\decoded_imm[30] ),
    .Y(_20677_));
 sky130_fd_sc_hd__clkbuf_2 _25648_ (.A(_20225_),
    .X(_20678_));
 sky130_fd_sc_hd__nor2_1 _25649_ (.A(_20678_),
    .B(_20477_),
    .Y(_20679_));
 sky130_fd_sc_hd__nor2_1 _25650_ (.A(_20677_),
    .B(_20679_),
    .Y(_20680_));
 sky130_fd_sc_hd__o22ai_4 _25651_ (.A1(_19788_),
    .A2(\decoded_imm[29] ),
    .B1(_20665_),
    .B2(_20673_),
    .Y(_20681_));
 sky130_fd_sc_hd__nand2_1 _25652_ (.A(_20681_),
    .B(_20671_),
    .Y(_20682_));
 sky130_fd_sc_hd__xor2_1 _25653_ (.A(_20680_),
    .B(_20682_),
    .X(_01461_));
 sky130_vsdinv _25654_ (.A(\reg_pc[31] ),
    .Y(_20683_));
 sky130_fd_sc_hd__nor2_2 _25655_ (.A(_19776_),
    .B(_20683_),
    .Y(_01462_));
 sky130_vsdinv _25656_ (.A(_18451_),
    .Y(_20684_));
 sky130_fd_sc_hd__nor2_1 _25657_ (.A(_20684_),
    .B(_20478_),
    .Y(_20685_));
 sky130_fd_sc_hd__nor2_1 _25658_ (.A(_18451_),
    .B(\decoded_imm[31] ),
    .Y(_20686_));
 sky130_fd_sc_hd__a22oi_1 _25659_ (.A1(_20678_),
    .A2(_20477_),
    .B1(_20681_),
    .B2(_20671_),
    .Y(_20687_));
 sky130_fd_sc_hd__o22ai_1 _25660_ (.A1(_20685_),
    .A2(_20686_),
    .B1(_20679_),
    .B2(_20687_),
    .Y(_20688_));
 sky130_fd_sc_hd__nor2_1 _25661_ (.A(_20686_),
    .B(_20685_),
    .Y(_20689_));
 sky130_fd_sc_hd__o2bb2ai_1 _25662_ (.A1_N(_20671_),
    .A2_N(_20681_),
    .B1(_19787_),
    .B2(\decoded_imm[30] ),
    .Y(_20690_));
 sky130_fd_sc_hd__o211ai_1 _25663_ (.A1(_20678_),
    .A2(_20477_),
    .B1(_20689_),
    .C1(_20690_),
    .Y(_20691_));
 sky130_fd_sc_hd__nand2_1 _25664_ (.A(_20688_),
    .B(_20691_),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_1 _25665_ (.A(_20364_),
    .B(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__and2_1 _25666_ (.A(_20364_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__buf_2 _25667_ (.A(_18526_),
    .X(_20692_));
 sky130_fd_sc_hd__a21oi_1 _25668_ (.A1(_20364_),
    .A2(_01473_),
    .B1(_20692_),
    .Y(_01474_));
 sky130_fd_sc_hd__and2_1 _25669_ (.A(_20364_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__clkbuf_2 _25670_ (.A(_20363_),
    .X(_20693_));
 sky130_fd_sc_hd__and2_1 _25671_ (.A(_20693_),
    .B(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__and2_1 _25672_ (.A(_20693_),
    .B(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__and2_1 _25673_ (.A(_20693_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__and2_1 _25674_ (.A(_20693_),
    .B(_01489_),
    .X(_01490_));
 sky130_fd_sc_hd__and2_1 _25675_ (.A(_20693_),
    .B(_01492_),
    .X(_01493_));
 sky130_fd_sc_hd__and2_1 _25676_ (.A(_20693_),
    .B(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__buf_1 _25677_ (.A(_20363_),
    .X(_20694_));
 sky130_fd_sc_hd__and2_1 _25678_ (.A(_20694_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__and2_1 _25679_ (.A(_20694_),
    .B(_01501_),
    .X(_01502_));
 sky130_fd_sc_hd__and2_1 _25680_ (.A(_20694_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__and2_1 _25681_ (.A(_20694_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__and2_1 _25682_ (.A(_20694_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__and2_1 _25683_ (.A(_20694_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__buf_1 _25684_ (.A(_20363_),
    .X(_20695_));
 sky130_fd_sc_hd__and2_1 _25685_ (.A(_20695_),
    .B(_01516_),
    .X(_01517_));
 sky130_fd_sc_hd__and2_1 _25686_ (.A(_20695_),
    .B(_01519_),
    .X(_01520_));
 sky130_fd_sc_hd__and2_1 _25687_ (.A(_20695_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__and2_1 _25688_ (.A(_20695_),
    .B(_01525_),
    .X(_01526_));
 sky130_fd_sc_hd__and2_1 _25689_ (.A(_20695_),
    .B(_01528_),
    .X(_01529_));
 sky130_fd_sc_hd__and2_1 _25690_ (.A(_20695_),
    .B(_01531_),
    .X(_01532_));
 sky130_fd_sc_hd__buf_1 _25691_ (.A(latched_branch),
    .X(_20696_));
 sky130_fd_sc_hd__and2_1 _25692_ (.A(_20696_),
    .B(_01534_),
    .X(_01535_));
 sky130_fd_sc_hd__and2_1 _25693_ (.A(_20696_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__and2_1 _25694_ (.A(_20696_),
    .B(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__and2_1 _25695_ (.A(_20696_),
    .B(_01543_),
    .X(_01544_));
 sky130_fd_sc_hd__and2_1 _25696_ (.A(_20696_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and2_1 _25697_ (.A(_20696_),
    .B(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__and2_1 _25698_ (.A(_20363_),
    .B(_01552_),
    .X(_01553_));
 sky130_fd_sc_hd__and2_1 _25699_ (.A(_20363_),
    .B(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__or2_1 _25700_ (.A(_02590_),
    .B(\decoded_imm_uj[1] ),
    .X(_20697_));
 sky130_fd_sc_hd__nand2_1 _25701_ (.A(_02590_),
    .B(\decoded_imm_uj[1] ),
    .Y(_20698_));
 sky130_fd_sc_hd__and2_1 _25702_ (.A(_20697_),
    .B(_20698_),
    .X(_01557_));
 sky130_fd_sc_hd__nor2_1 _25703_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .Y(_20699_));
 sky130_fd_sc_hd__and2_1 _25704_ (.A(_02560_),
    .B(\decoded_imm_uj[2] ),
    .X(_20700_));
 sky130_fd_sc_hd__nor2_2 _25705_ (.A(_20699_),
    .B(_20700_),
    .Y(_20701_));
 sky130_fd_sc_hd__xnor2_1 _25706_ (.A(_20698_),
    .B(_20701_),
    .Y(_01562_));
 sky130_fd_sc_hd__xor2_1 _25707_ (.A(_01561_),
    .B(_02410_),
    .X(_01565_));
 sky130_fd_sc_hd__nor2_1 _25708_ (.A(_02571_),
    .B(_02560_),
    .Y(_20702_));
 sky130_fd_sc_hd__nor2_1 _25709_ (.A(_18862_),
    .B(_01561_),
    .Y(_20703_));
 sky130_fd_sc_hd__nor2_1 _25710_ (.A(_20702_),
    .B(_20703_),
    .Y(_01567_));
 sky130_fd_sc_hd__xor2_1 _25711_ (.A(_02571_),
    .B(\decoded_imm_uj[3] ),
    .X(_20704_));
 sky130_fd_sc_hd__a31o_1 _25712_ (.A1(_20701_),
    .A2(_02590_),
    .A3(\decoded_imm_uj[1] ),
    .B1(_20700_),
    .X(_20705_));
 sky130_fd_sc_hd__xor2_1 _25713_ (.A(_20704_),
    .B(_20705_),
    .X(_01568_));
 sky130_fd_sc_hd__and3_1 _25714_ (.A(_02582_),
    .B(_02571_),
    .C(_02560_),
    .X(_20706_));
 sky130_fd_sc_hd__nor2_1 _25715_ (.A(_02582_),
    .B(_20703_),
    .Y(_20707_));
 sky130_fd_sc_hd__nor2_1 _25716_ (.A(_20706_),
    .B(_20707_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor2_2 _25717_ (.A(_01475_),
    .B(_00367_),
    .Y(_20708_));
 sky130_fd_sc_hd__nor2_1 _25718_ (.A(\decoded_imm_uj[4] ),
    .B(_02582_),
    .Y(_20709_));
 sky130_fd_sc_hd__or2_1 _25719_ (.A(_20708_),
    .B(_20709_),
    .X(_20710_));
 sky130_vsdinv _25720_ (.A(\decoded_imm_uj[3] ),
    .Y(_20711_));
 sky130_fd_sc_hd__o21ai_1 _25721_ (.A1(_02571_),
    .A2(\decoded_imm_uj[3] ),
    .B1(_20705_),
    .Y(_20712_));
 sky130_fd_sc_hd__o21a_1 _25722_ (.A1(_18862_),
    .A2(_20711_),
    .B1(_20712_),
    .X(_20713_));
 sky130_fd_sc_hd__xor2_1 _25723_ (.A(_20710_),
    .B(_20713_),
    .X(_01572_));
 sky130_fd_sc_hd__or2_1 _25724_ (.A(_02583_),
    .B(_20706_),
    .X(_20714_));
 sky130_fd_sc_hd__nand2_1 _25725_ (.A(_20706_),
    .B(_02583_),
    .Y(_20715_));
 sky130_fd_sc_hd__and2_1 _25726_ (.A(_20714_),
    .B(_20715_),
    .X(_01575_));
 sky130_fd_sc_hd__nor2_1 _25727_ (.A(_20709_),
    .B(_20713_),
    .Y(_20716_));
 sky130_fd_sc_hd__nor2_1 _25728_ (.A(_02583_),
    .B(\decoded_imm_uj[5] ),
    .Y(_20717_));
 sky130_fd_sc_hd__nand2_1 _25729_ (.A(_02583_),
    .B(\decoded_imm_uj[5] ),
    .Y(_20718_));
 sky130_fd_sc_hd__or2b_1 _25730_ (.A(_20717_),
    .B_N(_20718_),
    .X(_20719_));
 sky130_fd_sc_hd__o21ai_1 _25731_ (.A1(_20708_),
    .A2(_20716_),
    .B1(_20719_),
    .Y(_20720_));
 sky130_fd_sc_hd__or3_2 _25732_ (.A(_20708_),
    .B(_20719_),
    .C(_20716_),
    .X(_20721_));
 sky130_fd_sc_hd__nand2_1 _25733_ (.A(_20720_),
    .B(_20721_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _25734_ (.A(_18857_),
    .B(_20715_),
    .Y(_20722_));
 sky130_fd_sc_hd__and2_1 _25735_ (.A(_20715_),
    .B(_18857_),
    .X(_20723_));
 sky130_fd_sc_hd__nor2_1 _25736_ (.A(_20722_),
    .B(_20723_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_1 _25737_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .Y(_20724_));
 sky130_fd_sc_hd__and2_1 _25738_ (.A(_02584_),
    .B(\decoded_imm_uj[6] ),
    .X(_20725_));
 sky130_fd_sc_hd__nor2_1 _25739_ (.A(_20724_),
    .B(_20725_),
    .Y(_20726_));
 sky130_fd_sc_hd__o21bai_1 _25740_ (.A1(_20708_),
    .A2(_20716_),
    .B1_N(_20717_),
    .Y(_20727_));
 sky130_fd_sc_hd__nand2_1 _25741_ (.A(_20727_),
    .B(_20718_),
    .Y(_20728_));
 sky130_fd_sc_hd__xor2_1 _25742_ (.A(_20726_),
    .B(_20728_),
    .X(_01580_));
 sky130_fd_sc_hd__or2_1 _25743_ (.A(_02585_),
    .B(_20722_),
    .X(_20729_));
 sky130_fd_sc_hd__nand2_1 _25744_ (.A(_20722_),
    .B(_02585_),
    .Y(_20730_));
 sky130_fd_sc_hd__and2_1 _25745_ (.A(_20729_),
    .B(_20730_),
    .X(_01583_));
 sky130_fd_sc_hd__or2_1 _25746_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .X(_20731_));
 sky130_fd_sc_hd__nand2_2 _25747_ (.A(_02585_),
    .B(\decoded_imm_uj[7] ),
    .Y(_20732_));
 sky130_fd_sc_hd__nand2_1 _25748_ (.A(_20731_),
    .B(_20732_),
    .Y(_20733_));
 sky130_fd_sc_hd__a21oi_2 _25749_ (.A1(_20727_),
    .A2(_20718_),
    .B1(_20724_),
    .Y(_20734_));
 sky130_fd_sc_hd__nor2_1 _25750_ (.A(_20725_),
    .B(_20734_),
    .Y(_20735_));
 sky130_fd_sc_hd__xor2_1 _25751_ (.A(_20733_),
    .B(_20735_),
    .X(_01584_));
 sky130_fd_sc_hd__nor2_2 _25752_ (.A(_18852_),
    .B(_20730_),
    .Y(_20736_));
 sky130_fd_sc_hd__and2_1 _25753_ (.A(_20730_),
    .B(_18852_),
    .X(_20737_));
 sky130_fd_sc_hd__nor2_1 _25754_ (.A(_20736_),
    .B(_20737_),
    .Y(_01587_));
 sky130_fd_sc_hd__nor2_1 _25755_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .Y(_20738_));
 sky130_fd_sc_hd__and2_1 _25756_ (.A(_02586_),
    .B(\decoded_imm_uj[8] ),
    .X(_20739_));
 sky130_fd_sc_hd__nor2_1 _25757_ (.A(_20738_),
    .B(_20739_),
    .Y(_20740_));
 sky130_fd_sc_hd__o21ai_2 _25758_ (.A1(_20725_),
    .A2(_20734_),
    .B1(_20731_),
    .Y(_20741_));
 sky130_fd_sc_hd__nand2_1 _25759_ (.A(_20741_),
    .B(_20732_),
    .Y(_20742_));
 sky130_fd_sc_hd__xor2_1 _25760_ (.A(_20740_),
    .B(_20742_),
    .X(_01588_));
 sky130_fd_sc_hd__nor2_1 _25761_ (.A(_02587_),
    .B(_20736_),
    .Y(_20743_));
 sky130_fd_sc_hd__nand2_1 _25762_ (.A(_20736_),
    .B(_02587_),
    .Y(_20744_));
 sky130_vsdinv _25763_ (.A(_20744_),
    .Y(_20745_));
 sky130_fd_sc_hd__nor2_1 _25764_ (.A(_20743_),
    .B(_20745_),
    .Y(_01591_));
 sky130_fd_sc_hd__or2_1 _25765_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .X(_20746_));
 sky130_fd_sc_hd__nand2_2 _25766_ (.A(_02587_),
    .B(\decoded_imm_uj[9] ),
    .Y(_20747_));
 sky130_fd_sc_hd__nand2_1 _25767_ (.A(_20746_),
    .B(_20747_),
    .Y(_20748_));
 sky130_fd_sc_hd__a21oi_2 _25768_ (.A1(_20741_),
    .A2(_20732_),
    .B1(_20738_),
    .Y(_20749_));
 sky130_fd_sc_hd__nor2_1 _25769_ (.A(_20739_),
    .B(_20749_),
    .Y(_20750_));
 sky130_fd_sc_hd__xor2_1 _25770_ (.A(_20748_),
    .B(_20750_),
    .X(_01592_));
 sky130_fd_sc_hd__nor2_2 _25771_ (.A(_18848_),
    .B(_20744_),
    .Y(_20751_));
 sky130_fd_sc_hd__nor2_1 _25772_ (.A(_02588_),
    .B(_20745_),
    .Y(_20752_));
 sky130_fd_sc_hd__nor2_1 _25773_ (.A(_20751_),
    .B(_20752_),
    .Y(_01595_));
 sky130_fd_sc_hd__nor2_2 _25774_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .Y(_20753_));
 sky130_fd_sc_hd__and2_1 _25775_ (.A(_02588_),
    .B(\decoded_imm_uj[10] ),
    .X(_20754_));
 sky130_fd_sc_hd__nor2_1 _25776_ (.A(_20753_),
    .B(_20754_),
    .Y(_20755_));
 sky130_fd_sc_hd__o21ai_2 _25777_ (.A1(_20739_),
    .A2(_20749_),
    .B1(_20746_),
    .Y(_20756_));
 sky130_fd_sc_hd__nand2_1 _25778_ (.A(_20756_),
    .B(_20747_),
    .Y(_20757_));
 sky130_fd_sc_hd__xor2_1 _25779_ (.A(_20755_),
    .B(_20757_),
    .X(_01596_));
 sky130_fd_sc_hd__or2_1 _25780_ (.A(_02589_),
    .B(_20751_),
    .X(_20758_));
 sky130_fd_sc_hd__nand2_1 _25781_ (.A(_20751_),
    .B(_02589_),
    .Y(_20759_));
 sky130_fd_sc_hd__and2_1 _25782_ (.A(_20758_),
    .B(_20759_),
    .X(_01599_));
 sky130_vsdinv _25783_ (.A(\decoded_imm_uj[11] ),
    .Y(_20760_));
 sky130_fd_sc_hd__nor2_2 _25784_ (.A(_02589_),
    .B(_20760_),
    .Y(_20761_));
 sky130_fd_sc_hd__nor2_2 _25785_ (.A(\decoded_imm_uj[11] ),
    .B(_18846_),
    .Y(_20762_));
 sky130_fd_sc_hd__a21oi_4 _25786_ (.A1(_20756_),
    .A2(_20747_),
    .B1(_20753_),
    .Y(_20763_));
 sky130_fd_sc_hd__or4_1 _25787_ (.A(_20754_),
    .B(_20761_),
    .C(_20762_),
    .D(_20763_),
    .X(_20764_));
 sky130_fd_sc_hd__o22ai_4 _25788_ (.A1(_20761_),
    .A2(_20762_),
    .B1(_20754_),
    .B2(_20763_),
    .Y(_20765_));
 sky130_fd_sc_hd__and2_1 _25789_ (.A(_20764_),
    .B(_20765_),
    .X(_01600_));
 sky130_fd_sc_hd__nor2_2 _25790_ (.A(_18843_),
    .B(_20759_),
    .Y(_20766_));
 sky130_fd_sc_hd__and2_1 _25791_ (.A(_20759_),
    .B(_18843_),
    .X(_20767_));
 sky130_fd_sc_hd__nor2_1 _25792_ (.A(_20766_),
    .B(_20767_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _25793_ (.A(_18846_),
    .B(_20760_),
    .Y(_20768_));
 sky130_vsdinv _25794_ (.A(_20768_),
    .Y(_20769_));
 sky130_fd_sc_hd__nor2_1 _25795_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .Y(_20770_));
 sky130_fd_sc_hd__and2_1 _25796_ (.A(_02561_),
    .B(\decoded_imm_uj[12] ),
    .X(_20771_));
 sky130_fd_sc_hd__or2_2 _25797_ (.A(_20770_),
    .B(_20771_),
    .X(_20772_));
 sky130_fd_sc_hd__a21oi_4 _25798_ (.A1(_20765_),
    .A2(_20769_),
    .B1(_20772_),
    .Y(_20773_));
 sky130_fd_sc_hd__and3_1 _25799_ (.A(_20765_),
    .B(_20769_),
    .C(_20772_),
    .X(_20774_));
 sky130_fd_sc_hd__nor2_1 _25800_ (.A(_20773_),
    .B(_20774_),
    .Y(_01604_));
 sky130_fd_sc_hd__nor2_1 _25801_ (.A(_02562_),
    .B(_20766_),
    .Y(_20775_));
 sky130_fd_sc_hd__nand2_1 _25802_ (.A(_20766_),
    .B(_02562_),
    .Y(_20776_));
 sky130_vsdinv _25803_ (.A(_20776_),
    .Y(_20777_));
 sky130_fd_sc_hd__nor2_1 _25804_ (.A(_20775_),
    .B(_20777_),
    .Y(_01607_));
 sky130_vsdinv _25805_ (.A(\decoded_imm_uj[13] ),
    .Y(_20778_));
 sky130_fd_sc_hd__nor2_2 _25806_ (.A(_02562_),
    .B(_20778_),
    .Y(_20779_));
 sky130_fd_sc_hd__nor2_2 _25807_ (.A(\decoded_imm_uj[13] ),
    .B(_18841_),
    .Y(_20780_));
 sky130_fd_sc_hd__or4_1 _25808_ (.A(_20771_),
    .B(_20779_),
    .C(_20780_),
    .D(_20773_),
    .X(_20781_));
 sky130_fd_sc_hd__o22ai_4 _25809_ (.A1(_20779_),
    .A2(_20780_),
    .B1(_20771_),
    .B2(_20773_),
    .Y(_20782_));
 sky130_fd_sc_hd__and2_1 _25810_ (.A(_20781_),
    .B(_20782_),
    .X(_01608_));
 sky130_fd_sc_hd__nor2_2 _25811_ (.A(_18838_),
    .B(_20776_),
    .Y(_20783_));
 sky130_fd_sc_hd__nor2_1 _25812_ (.A(_02563_),
    .B(_20777_),
    .Y(_20784_));
 sky130_fd_sc_hd__nor2_1 _25813_ (.A(_20783_),
    .B(_20784_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2_1 _25814_ (.A(_18841_),
    .B(_20778_),
    .Y(_20785_));
 sky130_vsdinv _25815_ (.A(_20785_),
    .Y(_20786_));
 sky130_fd_sc_hd__nor2_1 _25816_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .Y(_20787_));
 sky130_fd_sc_hd__and2_1 _25817_ (.A(_02563_),
    .B(\decoded_imm_uj[14] ),
    .X(_20788_));
 sky130_fd_sc_hd__or2_2 _25818_ (.A(_20787_),
    .B(_20788_),
    .X(_20789_));
 sky130_fd_sc_hd__a21oi_4 _25819_ (.A1(_20782_),
    .A2(_20786_),
    .B1(_20789_),
    .Y(_20790_));
 sky130_fd_sc_hd__and3_1 _25820_ (.A(_20782_),
    .B(_20786_),
    .C(_20789_),
    .X(_20791_));
 sky130_fd_sc_hd__nor2_1 _25821_ (.A(_20790_),
    .B(_20791_),
    .Y(_01612_));
 sky130_fd_sc_hd__or2_1 _25822_ (.A(_02564_),
    .B(_20783_),
    .X(_20792_));
 sky130_fd_sc_hd__nand2_1 _25823_ (.A(_20783_),
    .B(_02564_),
    .Y(_20793_));
 sky130_fd_sc_hd__and2_1 _25824_ (.A(_20792_),
    .B(_20793_),
    .X(_01615_));
 sky130_fd_sc_hd__nor2_2 _25825_ (.A(_02564_),
    .B(_19715_),
    .Y(_20794_));
 sky130_fd_sc_hd__nor2_2 _25826_ (.A(\decoded_imm_uj[15] ),
    .B(_18835_),
    .Y(_20795_));
 sky130_fd_sc_hd__or4_4 _25827_ (.A(_20788_),
    .B(_20794_),
    .C(_20795_),
    .D(_20790_),
    .X(_20796_));
 sky130_fd_sc_hd__o22ai_4 _25828_ (.A1(_20794_),
    .A2(_20795_),
    .B1(_20788_),
    .B2(_20790_),
    .Y(_20797_));
 sky130_fd_sc_hd__and2_1 _25829_ (.A(_20796_),
    .B(_20797_),
    .X(_01616_));
 sky130_fd_sc_hd__nor2_2 _25830_ (.A(_18833_),
    .B(_20793_),
    .Y(_20798_));
 sky130_fd_sc_hd__and2_1 _25831_ (.A(_20793_),
    .B(_18833_),
    .X(_20799_));
 sky130_fd_sc_hd__nor2_1 _25832_ (.A(_20798_),
    .B(_20799_),
    .Y(_01619_));
 sky130_fd_sc_hd__nor2_1 _25833_ (.A(_18835_),
    .B(_19715_),
    .Y(_20800_));
 sky130_vsdinv _25834_ (.A(_20800_),
    .Y(_20801_));
 sky130_fd_sc_hd__nor2_1 _25835_ (.A(_02565_),
    .B(\decoded_imm_uj[16] ),
    .Y(_20802_));
 sky130_fd_sc_hd__nor2_4 _25836_ (.A(_18833_),
    .B(_19714_),
    .Y(_20803_));
 sky130_fd_sc_hd__nor2_1 _25837_ (.A(_20802_),
    .B(_20803_),
    .Y(_20804_));
 sky130_fd_sc_hd__a21boi_4 _25838_ (.A1(_20797_),
    .A2(_20801_),
    .B1_N(_20804_),
    .Y(_20805_));
 sky130_fd_sc_hd__o211a_1 _25839_ (.A1(_20803_),
    .A2(_20802_),
    .B1(_20801_),
    .C1(_20797_),
    .X(_20806_));
 sky130_fd_sc_hd__nor2_1 _25840_ (.A(_20805_),
    .B(_20806_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_1 _25841_ (.A(_02566_),
    .B(_20798_),
    .Y(_20807_));
 sky130_fd_sc_hd__nand2_1 _25842_ (.A(_20798_),
    .B(_02566_),
    .Y(_20808_));
 sky130_vsdinv _25843_ (.A(_20808_),
    .Y(_20809_));
 sky130_fd_sc_hd__nor2_1 _25844_ (.A(_20807_),
    .B(_20809_),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_2 _25845_ (.A(_02566_),
    .B(_19713_),
    .Y(_20810_));
 sky130_fd_sc_hd__nor2_2 _25846_ (.A(\decoded_imm_uj[17] ),
    .B(_18831_),
    .Y(_20811_));
 sky130_fd_sc_hd__or4_1 _25847_ (.A(_20803_),
    .B(_20810_),
    .C(_20811_),
    .D(_20805_),
    .X(_20812_));
 sky130_fd_sc_hd__o22ai_4 _25848_ (.A1(_20810_),
    .A2(_20811_),
    .B1(_20803_),
    .B2(_20805_),
    .Y(_20813_));
 sky130_fd_sc_hd__and2_1 _25849_ (.A(_20812_),
    .B(_20813_),
    .X(_01624_));
 sky130_fd_sc_hd__nor2_2 _25850_ (.A(_18828_),
    .B(_20808_),
    .Y(_20814_));
 sky130_fd_sc_hd__nor2_1 _25851_ (.A(_02567_),
    .B(_20809_),
    .Y(_20815_));
 sky130_fd_sc_hd__nor2_1 _25852_ (.A(_20814_),
    .B(_20815_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_1 _25853_ (.A(_02567_),
    .B(\decoded_imm_uj[18] ),
    .Y(_20816_));
 sky130_fd_sc_hd__nor2_4 _25854_ (.A(_18828_),
    .B(_19712_),
    .Y(_20817_));
 sky130_fd_sc_hd__nor2_1 _25855_ (.A(_20816_),
    .B(_20817_),
    .Y(_20818_));
 sky130_fd_sc_hd__nor2_1 _25856_ (.A(_18831_),
    .B(_19713_),
    .Y(_20819_));
 sky130_vsdinv _25857_ (.A(_20819_),
    .Y(_20820_));
 sky130_fd_sc_hd__nand2_1 _25858_ (.A(_20813_),
    .B(_20820_),
    .Y(_20821_));
 sky130_fd_sc_hd__xor2_1 _25859_ (.A(_20818_),
    .B(_20821_),
    .X(_01628_));
 sky130_fd_sc_hd__or2_1 _25860_ (.A(_02568_),
    .B(_20814_),
    .X(_20822_));
 sky130_fd_sc_hd__nand2_1 _25861_ (.A(_20814_),
    .B(_02568_),
    .Y(_20823_));
 sky130_fd_sc_hd__and2_1 _25862_ (.A(_20822_),
    .B(_20823_),
    .X(_01631_));
 sky130_vsdinv _25863_ (.A(\decoded_imm_uj[19] ),
    .Y(_20824_));
 sky130_fd_sc_hd__nor2_2 _25864_ (.A(_02568_),
    .B(_20824_),
    .Y(_20825_));
 sky130_fd_sc_hd__nor2_2 _25865_ (.A(\decoded_imm_uj[19] ),
    .B(_18826_),
    .Y(_20826_));
 sky130_fd_sc_hd__a22oi_4 _25866_ (.A1(_18828_),
    .A2(_19712_),
    .B1(_20813_),
    .B2(_20820_),
    .Y(_20827_));
 sky130_fd_sc_hd__or4_1 _25867_ (.A(_20817_),
    .B(_20825_),
    .C(_20826_),
    .D(_20827_),
    .X(_20828_));
 sky130_fd_sc_hd__o22ai_4 _25868_ (.A1(_20825_),
    .A2(_20826_),
    .B1(_20817_),
    .B2(_20827_),
    .Y(_20829_));
 sky130_fd_sc_hd__and2_1 _25869_ (.A(_20828_),
    .B(_20829_),
    .X(_01632_));
 sky130_fd_sc_hd__nor2_2 _25870_ (.A(_18823_),
    .B(_20823_),
    .Y(_20830_));
 sky130_fd_sc_hd__and2_1 _25871_ (.A(_20823_),
    .B(_18823_),
    .X(_20831_));
 sky130_fd_sc_hd__nor2_1 _25872_ (.A(_20830_),
    .B(_20831_),
    .Y(_01635_));
 sky130_fd_sc_hd__nor2_1 _25873_ (.A(_18826_),
    .B(_20824_),
    .Y(_20832_));
 sky130_vsdinv _25874_ (.A(_20832_),
    .Y(_20833_));
 sky130_fd_sc_hd__nor2_1 _25875_ (.A(_02569_),
    .B(_19711_),
    .Y(_20834_));
 sky130_fd_sc_hd__nor2_4 _25876_ (.A(_18823_),
    .B(_20079_),
    .Y(_20835_));
 sky130_fd_sc_hd__or2_1 _25877_ (.A(_20834_),
    .B(_20835_),
    .X(_20836_));
 sky130_fd_sc_hd__a21oi_1 _25878_ (.A1(_20829_),
    .A2(_20833_),
    .B1(_20836_),
    .Y(_20837_));
 sky130_fd_sc_hd__and3_1 _25879_ (.A(_20829_),
    .B(_20833_),
    .C(_20836_),
    .X(_20838_));
 sky130_fd_sc_hd__nor2_1 _25880_ (.A(_20837_),
    .B(_20838_),
    .Y(_01636_));
 sky130_fd_sc_hd__nor2_1 _25881_ (.A(_02570_),
    .B(_20830_),
    .Y(_20839_));
 sky130_fd_sc_hd__nand2_1 _25882_ (.A(_20830_),
    .B(_02570_),
    .Y(_20840_));
 sky130_vsdinv _25883_ (.A(_20840_),
    .Y(_20841_));
 sky130_fd_sc_hd__nor2_1 _25884_ (.A(_20839_),
    .B(_20841_),
    .Y(_01639_));
 sky130_fd_sc_hd__nor2_1 _25885_ (.A(_02570_),
    .B(_19709_),
    .Y(_20842_));
 sky130_fd_sc_hd__nor2_1 _25886_ (.A(_18820_),
    .B(_20078_),
    .Y(_20843_));
 sky130_fd_sc_hd__or2_1 _25887_ (.A(_20842_),
    .B(_20843_),
    .X(_20844_));
 sky130_vsdinv _25888_ (.A(_20844_),
    .Y(_20845_));
 sky130_fd_sc_hd__a22oi_4 _25889_ (.A1(_18823_),
    .A2(_20079_),
    .B1(_20829_),
    .B2(_20833_),
    .Y(_20846_));
 sky130_fd_sc_hd__or2_1 _25890_ (.A(_20835_),
    .B(_20846_),
    .X(_20847_));
 sky130_fd_sc_hd__or2_1 _25891_ (.A(_20845_),
    .B(_20847_),
    .X(_20848_));
 sky130_fd_sc_hd__nand2_1 _25892_ (.A(_20847_),
    .B(_20845_),
    .Y(_20849_));
 sky130_fd_sc_hd__and2_1 _25893_ (.A(_20848_),
    .B(_20849_),
    .X(_01640_));
 sky130_fd_sc_hd__nor2_1 _25894_ (.A(_18818_),
    .B(_20840_),
    .Y(_20850_));
 sky130_fd_sc_hd__nor2_1 _25895_ (.A(_02572_),
    .B(_20841_),
    .Y(_20851_));
 sky130_fd_sc_hd__nor2_1 _25896_ (.A(_20850_),
    .B(_20851_),
    .Y(_01643_));
 sky130_fd_sc_hd__xor2_4 _25897_ (.A(_02572_),
    .B(_19709_),
    .X(_20852_));
 sky130_vsdinv _25898_ (.A(_20852_),
    .Y(_20853_));
 sky130_fd_sc_hd__a21oi_1 _25899_ (.A1(_20847_),
    .A2(_20845_),
    .B1(_20843_),
    .Y(_20854_));
 sky130_fd_sc_hd__xor2_1 _25900_ (.A(_20853_),
    .B(_20854_),
    .X(_01644_));
 sky130_fd_sc_hd__or2_1 _25901_ (.A(_02573_),
    .B(_20850_),
    .X(_20855_));
 sky130_fd_sc_hd__nand2_1 _25902_ (.A(_20850_),
    .B(_02573_),
    .Y(_20856_));
 sky130_fd_sc_hd__and2_1 _25903_ (.A(_20855_),
    .B(_20856_),
    .X(_01647_));
 sky130_fd_sc_hd__nor2_2 _25904_ (.A(_18816_),
    .B(_20078_),
    .Y(_20857_));
 sky130_vsdinv _25905_ (.A(_20857_),
    .Y(_20858_));
 sky130_fd_sc_hd__nand2_1 _25906_ (.A(_18816_),
    .B(_20078_),
    .Y(_20859_));
 sky130_fd_sc_hd__nand2_1 _25907_ (.A(_20858_),
    .B(_20859_),
    .Y(_20860_));
 sky130_vsdinv _25908_ (.A(_20860_),
    .Y(_20861_));
 sky130_fd_sc_hd__o21a_1 _25909_ (.A1(_02572_),
    .A2(_02570_),
    .B1(_19710_),
    .X(_20862_));
 sky130_fd_sc_hd__nor2_1 _25910_ (.A(_20853_),
    .B(_20849_),
    .Y(_20863_));
 sky130_fd_sc_hd__nor3_1 _25911_ (.A(_20861_),
    .B(_20862_),
    .C(_20863_),
    .Y(_20864_));
 sky130_fd_sc_hd__o21a_1 _25912_ (.A1(_20862_),
    .A2(_20863_),
    .B1(_20861_),
    .X(_20865_));
 sky130_fd_sc_hd__nor2_1 _25913_ (.A(_20864_),
    .B(_20865_),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_2 _25914_ (.A(_18813_),
    .B(_20856_),
    .Y(_20866_));
 sky130_fd_sc_hd__and2_1 _25915_ (.A(_20856_),
    .B(_18813_),
    .X(_20867_));
 sky130_fd_sc_hd__nor2_1 _25916_ (.A(_20866_),
    .B(_20867_),
    .Y(_01651_));
 sky130_fd_sc_hd__xor2_2 _25917_ (.A(_02574_),
    .B(_19709_),
    .X(_20868_));
 sky130_fd_sc_hd__nor3_1 _25918_ (.A(_20857_),
    .B(_20868_),
    .C(_20865_),
    .Y(_20869_));
 sky130_fd_sc_hd__o21a_1 _25919_ (.A1(_20857_),
    .A2(_20865_),
    .B1(_20868_),
    .X(_20870_));
 sky130_fd_sc_hd__nor2_1 _25920_ (.A(_20869_),
    .B(_20870_),
    .Y(_01652_));
 sky130_fd_sc_hd__nor2_1 _25921_ (.A(_02575_),
    .B(_20866_),
    .Y(_20871_));
 sky130_fd_sc_hd__nand2_1 _25922_ (.A(_20866_),
    .B(_02575_),
    .Y(_20872_));
 sky130_vsdinv _25923_ (.A(_20872_),
    .Y(_20873_));
 sky130_fd_sc_hd__nor2_1 _25924_ (.A(_20871_),
    .B(_20873_),
    .Y(_01655_));
 sky130_fd_sc_hd__nor2_2 _25925_ (.A(_02575_),
    .B(_20079_),
    .Y(_20874_));
 sky130_fd_sc_hd__nor2_2 _25926_ (.A(_19710_),
    .B(_18811_),
    .Y(_20875_));
 sky130_fd_sc_hd__or2_1 _25927_ (.A(_20874_),
    .B(_20875_),
    .X(_20876_));
 sky130_fd_sc_hd__and3_1 _25928_ (.A(_20858_),
    .B(_20868_),
    .C(_20859_),
    .X(_20877_));
 sky130_fd_sc_hd__o2111ai_4 _25929_ (.A1(_20835_),
    .A2(_20846_),
    .B1(_20845_),
    .C1(_20852_),
    .D1(_20877_),
    .Y(_20878_));
 sky130_fd_sc_hd__a41o_1 _25930_ (.A1(_18813_),
    .A2(_18816_),
    .A3(_18818_),
    .A4(_18820_),
    .B1(_20079_),
    .X(_20879_));
 sky130_fd_sc_hd__nand2_2 _25931_ (.A(_20878_),
    .B(_20879_),
    .Y(_20880_));
 sky130_fd_sc_hd__or2_1 _25932_ (.A(_20876_),
    .B(_20880_),
    .X(_20881_));
 sky130_fd_sc_hd__nand2_1 _25933_ (.A(_20880_),
    .B(_20876_),
    .Y(_20882_));
 sky130_fd_sc_hd__and2_1 _25934_ (.A(_20881_),
    .B(_20882_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_2 _25935_ (.A(_18808_),
    .B(_20872_),
    .Y(_20883_));
 sky130_fd_sc_hd__nor2_1 _25936_ (.A(_02576_),
    .B(_20873_),
    .Y(_20884_));
 sky130_fd_sc_hd__nor2_1 _25937_ (.A(_20883_),
    .B(_20884_),
    .Y(_01659_));
 sky130_fd_sc_hd__xor2_4 _25938_ (.A(_02576_),
    .B(_19710_),
    .X(_20885_));
 sky130_fd_sc_hd__o21ai_1 _25939_ (.A1(_18811_),
    .A2(_20080_),
    .B1(_20882_),
    .Y(_20886_));
 sky130_fd_sc_hd__xor2_1 _25940_ (.A(_20885_),
    .B(_20886_),
    .X(_01660_));
 sky130_fd_sc_hd__or2_1 _25941_ (.A(_02577_),
    .B(_20883_),
    .X(_20887_));
 sky130_fd_sc_hd__nand2_1 _25942_ (.A(_20883_),
    .B(_02577_),
    .Y(_20888_));
 sky130_fd_sc_hd__and2_1 _25943_ (.A(_20887_),
    .B(_20888_),
    .X(_01663_));
 sky130_fd_sc_hd__nand3_2 _25944_ (.A(_20880_),
    .B(_20876_),
    .C(_20885_),
    .Y(_20889_));
 sky130_fd_sc_hd__o21a_1 _25945_ (.A1(_02576_),
    .A2(_02575_),
    .B1(_19710_),
    .X(_04073_));
 sky130_vsdinv _25946_ (.A(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__nor2_1 _25947_ (.A(_02577_),
    .B(_19709_),
    .Y(_04075_));
 sky130_fd_sc_hd__nor2_2 _25948_ (.A(_18805_),
    .B(_20079_),
    .Y(_04076_));
 sky130_fd_sc_hd__or2_1 _25949_ (.A(_04075_),
    .B(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__a21oi_2 _25950_ (.A1(_20889_),
    .A2(_04074_),
    .B1(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__and3_1 _25951_ (.A(_20889_),
    .B(_04077_),
    .C(_04074_),
    .X(_04079_));
 sky130_fd_sc_hd__nor2_1 _25952_ (.A(_04078_),
    .B(_04079_),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_1 _25953_ (.A(_18803_),
    .B(_20888_),
    .Y(_04080_));
 sky130_fd_sc_hd__and2_1 _25954_ (.A(_20888_),
    .B(_18803_),
    .X(_04081_));
 sky130_fd_sc_hd__nor2_1 _25955_ (.A(_04080_),
    .B(_04081_),
    .Y(_01667_));
 sky130_fd_sc_hd__xor2_2 _25956_ (.A(_02578_),
    .B(_19709_),
    .X(_04082_));
 sky130_fd_sc_hd__nor3_1 _25957_ (.A(_04076_),
    .B(_04082_),
    .C(_04078_),
    .Y(_04083_));
 sky130_fd_sc_hd__o21a_1 _25958_ (.A1(_04076_),
    .A2(_04078_),
    .B1(_04082_),
    .X(_04084_));
 sky130_fd_sc_hd__nor2_1 _25959_ (.A(_04083_),
    .B(_04084_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_1 _25960_ (.A(_02579_),
    .B(_04080_),
    .Y(_04085_));
 sky130_fd_sc_hd__and2_1 _25961_ (.A(_04080_),
    .B(_02579_),
    .X(_04086_));
 sky130_fd_sc_hd__nor2_1 _25962_ (.A(_04085_),
    .B(_04086_),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2_1 _25963_ (.A(_18801_),
    .B(_20080_),
    .Y(_04087_));
 sky130_fd_sc_hd__nand2_1 _25964_ (.A(_02579_),
    .B(_19710_),
    .Y(_04088_));
 sky130_fd_sc_hd__and2_1 _25965_ (.A(_04087_),
    .B(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__and2b_1 _25966_ (.A_N(_04077_),
    .B(_04082_),
    .X(_04090_));
 sky130_fd_sc_hd__o2111ai_4 _25967_ (.A1(_20874_),
    .A2(_20875_),
    .B1(_20885_),
    .C1(_04090_),
    .D1(_20880_),
    .Y(_04091_));
 sky130_fd_sc_hd__a41o_1 _25968_ (.A1(_18803_),
    .A2(_18805_),
    .A3(_18808_),
    .A4(_18811_),
    .B1(_20080_),
    .X(_04092_));
 sky130_fd_sc_hd__nand2_2 _25969_ (.A(_04091_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__or2_1 _25970_ (.A(_04089_),
    .B(_04093_),
    .X(_04094_));
 sky130_fd_sc_hd__nand2_1 _25971_ (.A(_04093_),
    .B(_04089_),
    .Y(_04095_));
 sky130_fd_sc_hd__and2_1 _25972_ (.A(_04094_),
    .B(_04095_),
    .X(_01672_));
 sky130_fd_sc_hd__or2_1 _25973_ (.A(_02580_),
    .B(_04086_),
    .X(_04096_));
 sky130_fd_sc_hd__nand2_1 _25974_ (.A(_04086_),
    .B(_02580_),
    .Y(_04097_));
 sky130_fd_sc_hd__and2_1 _25975_ (.A(_04096_),
    .B(_04097_),
    .X(_01675_));
 sky130_fd_sc_hd__nor2_1 _25976_ (.A(_02580_),
    .B(_19711_),
    .Y(_04098_));
 sky130_fd_sc_hd__nor2_1 _25977_ (.A(_18798_),
    .B(_20080_),
    .Y(_04099_));
 sky130_fd_sc_hd__nor2_1 _25978_ (.A(_04098_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__a21o_1 _25979_ (.A1(_04095_),
    .A2(_04088_),
    .B1(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__nand3_1 _25980_ (.A(_04095_),
    .B(_04088_),
    .C(_04100_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand2_1 _25981_ (.A(_04101_),
    .B(_04102_),
    .Y(_01676_));
 sky130_fd_sc_hd__xor2_1 _25982_ (.A(_18795_),
    .B(_04097_),
    .X(_01679_));
 sky130_fd_sc_hd__nand2_1 _25983_ (.A(_20080_),
    .B(_02581_),
    .Y(_04103_));
 sky130_fd_sc_hd__nand2_1 _25984_ (.A(_18795_),
    .B(_19711_),
    .Y(_04104_));
 sky130_vsdinv _25985_ (.A(_04098_),
    .Y(_04105_));
 sky130_fd_sc_hd__nand3_1 _25986_ (.A(_04093_),
    .B(_04089_),
    .C(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__o21a_1 _25987_ (.A1(_02580_),
    .A2(_02579_),
    .B1(_19711_),
    .X(_04107_));
 sky130_vsdinv _25988_ (.A(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__a22oi_1 _25989_ (.A1(_04103_),
    .A2(_04104_),
    .B1(_04106_),
    .B2(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__nand2_1 _25990_ (.A(_04103_),
    .B(_04104_),
    .Y(_04110_));
 sky130_fd_sc_hd__a311oi_4 _25991_ (.A1(_04093_),
    .A2(_04089_),
    .A3(_04105_),
    .B1(_04107_),
    .C1(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__nor2_1 _25992_ (.A(_04109_),
    .B(_04111_),
    .Y(_01680_));
 sky130_fd_sc_hd__buf_4 _25993_ (.A(\mem_wordsize[2] ),
    .X(_04112_));
 sky130_fd_sc_hd__nor2_4 _25994_ (.A(_04112_),
    .B(\mem_wordsize[1] ),
    .Y(_04113_));
 sky130_fd_sc_hd__clkbuf_4 _25995_ (.A(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__buf_4 _25996_ (.A(_04114_),
    .X(_01683_));
 sky130_fd_sc_hd__a21oi_4 _25997_ (.A1(_20338_),
    .A2(_04112_),
    .B1(_04113_),
    .Y(_04115_));
 sky130_fd_sc_hd__o21a_4 _25998_ (.A1(_19819_),
    .A2(_19820_),
    .B1(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__nor2_1 _25999_ (.A(_04116_),
    .B(_19473_),
    .Y(_01684_));
 sky130_fd_sc_hd__and3_1 _26000_ (.A(_00301_),
    .B(_20360_),
    .C(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__nor2_2 _26001_ (.A(_19819_),
    .B(_20119_),
    .Y(_04117_));
 sky130_vsdinv _26002_ (.A(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__nand2_8 _26003_ (.A(_04118_),
    .B(_04115_),
    .Y(net234));
 sky130_fd_sc_hd__and3_1 _26004_ (.A(net234),
    .B(_18630_),
    .C(_19472_),
    .X(_01687_));
 sky130_fd_sc_hd__and3_1 _26005_ (.A(_00301_),
    .B(_20360_),
    .C(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__nor2_2 _26006_ (.A(_19820_),
    .B(_20338_),
    .Y(_04119_));
 sky130_fd_sc_hd__nor2_1 _26007_ (.A(_20338_),
    .B(_20132_),
    .Y(_04120_));
 sky130_fd_sc_hd__or3_4 _26008_ (.A(_04113_),
    .B(_04119_),
    .C(_04120_),
    .X(net235));
 sky130_fd_sc_hd__and3_1 _26009_ (.A(net235),
    .B(_18630_),
    .C(_19472_),
    .X(_01690_));
 sky130_fd_sc_hd__and3_1 _26010_ (.A(_00301_),
    .B(_20360_),
    .C(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__nor2_2 _26011_ (.A(_20338_),
    .B(_20119_),
    .Y(_04121_));
 sky130_fd_sc_hd__or3_4 _26012_ (.A(_04114_),
    .B(_04120_),
    .C(_04121_),
    .X(net236));
 sky130_fd_sc_hd__and2_1 _26013_ (.A(net232),
    .B(net236),
    .X(_01693_));
 sky130_fd_sc_hd__and3_1 _26014_ (.A(_00301_),
    .B(_20360_),
    .C(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__nor2_4 _26015_ (.A(\irq_pending[1] ),
    .B(net12),
    .Y(_01696_));
 sky130_fd_sc_hd__inv_2 _26016_ (.A(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__nor2_1 _26017_ (.A(_18625_),
    .B(_01696_),
    .Y(_01698_));
 sky130_fd_sc_hd__clkbuf_4 _26018_ (.A(_20150_),
    .X(_04122_));
 sky130_fd_sc_hd__or3_4 _26019_ (.A(\cpu_state[0] ),
    .B(_02542_),
    .C(_18553_),
    .X(_04123_));
 sky130_fd_sc_hd__nor2_1 _26020_ (.A(_04122_),
    .B(_04123_),
    .Y(_01700_));
 sky130_fd_sc_hd__and2_1 _26021_ (.A(_20128_),
    .B(_01696_),
    .X(_01701_));
 sky130_fd_sc_hd__a2bb2o_1 _26022_ (.A1_N(_18520_),
    .A2_N(_01704_),
    .B1(_01697_),
    .B2(_04123_),
    .X(_01705_));
 sky130_vsdinv _26023_ (.A(net33),
    .Y(_01707_));
 sky130_fd_sc_hd__clkbuf_2 _26024_ (.A(_04121_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_2 _26025_ (.A(_04117_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_2 _26026_ (.A(_04119_),
    .X(_04126_));
 sky130_fd_sc_hd__a22o_1 _26027_ (.A1(_04125_),
    .A2(net63),
    .B1(net40),
    .B2(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__a21oi_1 _26028_ (.A1(net49),
    .A2(_04124_),
    .B1(_04127_),
    .Y(_01708_));
 sky130_fd_sc_hd__clkbuf_2 _26029_ (.A(_04112_),
    .X(_04128_));
 sky130_fd_sc_hd__o2bb2a_1 _26030_ (.A1_N(_04128_),
    .A2_N(_01710_),
    .B1(_01709_),
    .B2(_20359_),
    .X(_01711_));
 sky130_vsdinv _26031_ (.A(instr_rdinstrh),
    .Y(_04129_));
 sky130_fd_sc_hd__buf_2 _26032_ (.A(_04129_),
    .X(_04130_));
 sky130_vsdinv _26033_ (.A(_19760_),
    .Y(_04131_));
 sky130_fd_sc_hd__buf_2 _26034_ (.A(_04131_),
    .X(_04132_));
 sky130_vsdinv _26035_ (.A(instr_rdcycleh),
    .Y(_04133_));
 sky130_fd_sc_hd__clkbuf_2 _26036_ (.A(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__and3_4 _26037_ (.A(_04130_),
    .B(_04132_),
    .C(_04134_),
    .X(_01714_));
 sky130_fd_sc_hd__buf_2 _26038_ (.A(_04131_),
    .X(_04135_));
 sky130_fd_sc_hd__nand2_1 _26039_ (.A(\count_instr[32] ),
    .B(_19752_),
    .Y(_04136_));
 sky130_fd_sc_hd__o221a_1 _26040_ (.A1(_19055_),
    .A2(_04135_),
    .B1(_04134_),
    .B2(_19303_),
    .C1(_04136_),
    .X(_01715_));
 sky130_fd_sc_hd__nand2_1 _26041_ (.A(\irq_mask[0] ),
    .B(_19739_),
    .Y(_04137_));
 sky130_fd_sc_hd__o221a_1 _26042_ (.A1(_18492_),
    .A2(_20368_),
    .B1(_18489_),
    .B2(_18628_),
    .C1(_04137_),
    .X(_01718_));
 sky130_fd_sc_hd__clkbuf_4 _26043_ (.A(_18478_),
    .X(_04138_));
 sky130_fd_sc_hd__nand2_1 _26044_ (.A(\decoded_imm[0] ),
    .B(\reg_next_pc[0] ),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_1 _26045_ (.A(_20481_),
    .B(_20480_),
    .Y(_04140_));
 sky130_fd_sc_hd__buf_2 _26046_ (.A(_20150_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_4 _26047_ (.A(_18542_),
    .X(_04142_));
 sky130_fd_sc_hd__nor2_1 _26048_ (.A(_01719_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__clkbuf_4 _26049_ (.A(_18328_),
    .X(_04144_));
 sky130_fd_sc_hd__nor2_1 _26050_ (.A(_01712_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__a211o_1 _26051_ (.A1(_04141_),
    .A2(_01713_),
    .B1(_04143_),
    .C1(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__a31o_1 _26052_ (.A1(_04138_),
    .A2(_04139_),
    .A3(_04140_),
    .B1(_04146_),
    .X(_01720_));
 sky130_vsdinv _26053_ (.A(net44),
    .Y(_01721_));
 sky130_fd_sc_hd__a22o_1 _26054_ (.A1(_04125_),
    .A2(net64),
    .B1(net41),
    .B2(_04126_),
    .X(_04147_));
 sky130_fd_sc_hd__a21oi_1 _26055_ (.A1(net50),
    .A2(_04124_),
    .B1(_04147_),
    .Y(_01722_));
 sky130_fd_sc_hd__o2bb2a_1 _26056_ (.A1_N(_04128_),
    .A2_N(_01724_),
    .B1(_01723_),
    .B2(_20359_),
    .X(_01725_));
 sky130_fd_sc_hd__nand2_1 _26057_ (.A(\count_instr[33] ),
    .B(_19752_),
    .Y(_04148_));
 sky130_fd_sc_hd__o221a_1 _26058_ (.A1(_19081_),
    .A2(_04135_),
    .B1(_04134_),
    .B2(_19207_),
    .C1(_04148_),
    .X(_01729_));
 sky130_fd_sc_hd__clkbuf_2 _26059_ (.A(_18494_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_2 _26060_ (.A(_18492_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_2 _26061_ (.A(_18490_),
    .X(_04151_));
 sky130_fd_sc_hd__buf_2 _26062_ (.A(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__nand2_1 _26063_ (.A(\cpuregs_rs1[1] ),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__o221a_1 _26064_ (.A1(_18625_),
    .A2(_04149_),
    .B1(_04150_),
    .B2(_20367_),
    .C1(_04153_),
    .X(_01731_));
 sky130_fd_sc_hd__nor2_1 _26065_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_04154_));
 sky130_fd_sc_hd__nand2_1 _26066_ (.A(\reg_pc[1] ),
    .B(\decoded_imm[1] ),
    .Y(_04155_));
 sky130_fd_sc_hd__or2b_1 _26067_ (.A(_04154_),
    .B_N(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__or2_1 _26068_ (.A(_04139_),
    .B(_04156_),
    .X(_04157_));
 sky130_fd_sc_hd__buf_2 _26069_ (.A(_18478_),
    .X(_04158_));
 sky130_fd_sc_hd__nand2_1 _26070_ (.A(_04156_),
    .B(_04139_),
    .Y(_04159_));
 sky130_fd_sc_hd__clkbuf_4 _26071_ (.A(_19090_),
    .X(_04160_));
 sky130_fd_sc_hd__nor2_1 _26072_ (.A(_01732_),
    .B(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__clkbuf_4 _26073_ (.A(_18519_),
    .X(_04162_));
 sky130_fd_sc_hd__a2bb2o_1 _26074_ (.A1_N(_01726_),
    .A2_N(_20183_),
    .B1(_04162_),
    .B2(_01727_),
    .X(_04163_));
 sky130_fd_sc_hd__a311o_1 _26075_ (.A1(_04157_),
    .A2(_04158_),
    .A3(_04159_),
    .B1(_04161_),
    .C1(_04163_),
    .X(_01733_));
 sky130_vsdinv _26076_ (.A(net55),
    .Y(_01734_));
 sky130_fd_sc_hd__a22o_1 _26077_ (.A1(_04125_),
    .A2(net34),
    .B1(net42),
    .B2(_04126_),
    .X(_04164_));
 sky130_fd_sc_hd__a21oi_1 _26078_ (.A1(net51),
    .A2(_04124_),
    .B1(_04164_),
    .Y(_01735_));
 sky130_fd_sc_hd__o2bb2a_1 _26079_ (.A1_N(_04128_),
    .A2_N(_01737_),
    .B1(_01736_),
    .B2(_20359_),
    .X(_01738_));
 sky130_fd_sc_hd__nand2_1 _26080_ (.A(\count_instr[2] ),
    .B(_19761_),
    .Y(_04165_));
 sky130_fd_sc_hd__o221a_1 _26081_ (.A1(_18909_),
    .A2(_04130_),
    .B1(_04134_),
    .B2(_19208_),
    .C1(_04165_),
    .X(_01742_));
 sky130_fd_sc_hd__nand2_1 _26082_ (.A(\cpuregs_rs1[2] ),
    .B(_04152_),
    .Y(_04166_));
 sky130_fd_sc_hd__o221a_1 _26083_ (.A1(_18623_),
    .A2(_04149_),
    .B1(_04150_),
    .B2(_20405_),
    .C1(_04166_),
    .X(_01744_));
 sky130_fd_sc_hd__o21ai_1 _26084_ (.A1(_04139_),
    .A2(_04154_),
    .B1(_04155_),
    .Y(_04167_));
 sky130_fd_sc_hd__xor2_1 _26085_ (.A(\reg_pc[2] ),
    .B(\decoded_imm[2] ),
    .X(_04168_));
 sky130_fd_sc_hd__or2_1 _26086_ (.A(_04167_),
    .B(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__nand2_1 _26087_ (.A(_04168_),
    .B(_04167_),
    .Y(_04170_));
 sky130_fd_sc_hd__buf_2 _26088_ (.A(_18478_),
    .X(_04171_));
 sky130_fd_sc_hd__nor2_2 _26089_ (.A(_01745_),
    .B(_04160_),
    .Y(_04172_));
 sky130_fd_sc_hd__a2bb2o_1 _26090_ (.A1_N(_01739_),
    .A2_N(_20183_),
    .B1(_04162_),
    .B2(_01740_),
    .X(_04173_));
 sky130_fd_sc_hd__a311o_1 _26091_ (.A1(_04169_),
    .A2(_04170_),
    .A3(_04171_),
    .B1(_04172_),
    .C1(_04173_),
    .X(_01746_));
 sky130_vsdinv _26092_ (.A(net58),
    .Y(_01747_));
 sky130_fd_sc_hd__a22o_1 _26093_ (.A1(_04125_),
    .A2(net35),
    .B1(net515),
    .B2(_04126_),
    .X(_04174_));
 sky130_fd_sc_hd__a21oi_1 _26094_ (.A1(net52),
    .A2(_04124_),
    .B1(_04174_),
    .Y(_01748_));
 sky130_fd_sc_hd__o2bb2a_1 _26095_ (.A1_N(_04128_),
    .A2_N(_01750_),
    .B1(_01749_),
    .B2(_20359_),
    .X(_01751_));
 sky130_fd_sc_hd__buf_2 _26096_ (.A(_04131_),
    .X(_04175_));
 sky130_fd_sc_hd__nand2_1 _26097_ (.A(\count_instr[35] ),
    .B(_19752_),
    .Y(_04176_));
 sky130_fd_sc_hd__o221a_1 _26098_ (.A1(_19079_),
    .A2(_04175_),
    .B1(_04134_),
    .B2(_19297_),
    .C1(_04176_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _26099_ (.A(\cpuregs_rs1[3] ),
    .B(_04152_),
    .Y(_04177_));
 sky130_fd_sc_hd__o221a_1 _26100_ (.A1(_18418_),
    .A2(_04149_),
    .B1(_04150_),
    .B2(_20406_),
    .C1(_04177_),
    .X(_01757_));
 sky130_fd_sc_hd__nor2_1 _26101_ (.A(_01758_),
    .B(_04160_),
    .Y(_04178_));
 sky130_fd_sc_hd__nor2_1 _26102_ (.A(_01752_),
    .B(_20348_),
    .Y(_04179_));
 sky130_fd_sc_hd__nor2_2 _26103_ (.A(_20489_),
    .B(_20036_),
    .Y(_04180_));
 sky130_fd_sc_hd__o21ai_1 _26104_ (.A1(\reg_pc[2] ),
    .A2(\decoded_imm[2] ),
    .B1(_04167_),
    .Y(_04181_));
 sky130_fd_sc_hd__o21a_1 _26105_ (.A1(_02073_),
    .A2(_20029_),
    .B1(_04181_),
    .X(_04182_));
 sky130_fd_sc_hd__a21o_1 _26106_ (.A1(_20489_),
    .A2(_20036_),
    .B1(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__nor2_1 _26107_ (.A(\reg_pc[3] ),
    .B(\decoded_imm[3] ),
    .Y(_04184_));
 sky130_fd_sc_hd__o21ai_1 _26108_ (.A1(_04180_),
    .A2(_04184_),
    .B1(_04182_),
    .Y(_04185_));
 sky130_fd_sc_hd__o211a_1 _26109_ (.A1(_04180_),
    .A2(_04183_),
    .B1(_18478_),
    .C1(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__a2111o_1 _26110_ (.A1(_04122_),
    .A2(_01753_),
    .B1(_04178_),
    .C1(_04179_),
    .D1(_04186_),
    .X(_01759_));
 sky130_vsdinv _26111_ (.A(net59),
    .Y(_01760_));
 sky130_fd_sc_hd__a22o_1 _26112_ (.A1(_04125_),
    .A2(net517),
    .B1(net514),
    .B2(_04126_),
    .X(_04187_));
 sky130_fd_sc_hd__a21oi_1 _26113_ (.A1(net53),
    .A2(_04124_),
    .B1(_04187_),
    .Y(_01761_));
 sky130_fd_sc_hd__buf_2 _26114_ (.A(_04112_),
    .X(_04188_));
 sky130_fd_sc_hd__o2bb2a_1 _26115_ (.A1_N(_04188_),
    .A2_N(_01763_),
    .B1(_01762_),
    .B2(_20359_),
    .X(_01764_));
 sky130_fd_sc_hd__nand2_1 _26116_ (.A(\count_instr[36] ),
    .B(_19752_),
    .Y(_04189_));
 sky130_fd_sc_hd__o221a_1 _26117_ (.A1(_19054_),
    .A2(_04175_),
    .B1(_04134_),
    .B2(_19300_),
    .C1(_04189_),
    .X(_01768_));
 sky130_fd_sc_hd__clkbuf_4 _26118_ (.A(_04151_),
    .X(_04190_));
 sky130_fd_sc_hd__a22o_1 _26119_ (.A1(\irq_mask[4] ),
    .A2(_19739_),
    .B1(_19725_),
    .B2(\timer[4] ),
    .X(_04191_));
 sky130_fd_sc_hd__a21oi_1 _26120_ (.A1(\cpuregs_rs1[4] ),
    .A2(_04190_),
    .B1(_04191_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_1 _26121_ (.A(_20495_),
    .B(_20041_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand2_1 _26122_ (.A(\reg_pc[4] ),
    .B(\decoded_imm[4] ),
    .Y(_04193_));
 sky130_fd_sc_hd__nand2_1 _26123_ (.A(_04192_),
    .B(_04193_),
    .Y(_04194_));
 sky130_vsdinv _26124_ (.A(_04194_),
    .Y(_04195_));
 sky130_vsdinv _26125_ (.A(_04180_),
    .Y(_04196_));
 sky130_fd_sc_hd__nand2_2 _26126_ (.A(_04183_),
    .B(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__nor2_1 _26127_ (.A(_04195_),
    .B(_04197_),
    .Y(_04198_));
 sky130_vsdinv _26128_ (.A(_04197_),
    .Y(_04199_));
 sky130_fd_sc_hd__nor2_1 _26129_ (.A(_04194_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _26130_ (.A(_04141_),
    .B(_01766_),
    .Y(_04201_));
 sky130_fd_sc_hd__o221a_1 _26131_ (.A1(_01765_),
    .A2(_04144_),
    .B1(_19131_),
    .B2(_01771_),
    .C1(_04201_),
    .X(_04202_));
 sky130_fd_sc_hd__o31ai_2 _26132_ (.A1(_20195_),
    .A2(_04198_),
    .A3(_04200_),
    .B1(_04202_),
    .Y(_01772_));
 sky130_vsdinv _26133_ (.A(net512),
    .Y(_01773_));
 sky130_fd_sc_hd__a22o_1 _26134_ (.A1(_04125_),
    .A2(net37),
    .B1(net46),
    .B2(_04126_),
    .X(_04203_));
 sky130_fd_sc_hd__a21oi_1 _26135_ (.A1(net54),
    .A2(_04124_),
    .B1(_04203_),
    .Y(_01774_));
 sky130_fd_sc_hd__o2bb2a_1 _26136_ (.A1_N(_04188_),
    .A2_N(_01776_),
    .B1(_01775_),
    .B2(_20358_),
    .X(_01777_));
 sky130_fd_sc_hd__clkbuf_2 _26137_ (.A(_04133_),
    .X(_04204_));
 sky130_fd_sc_hd__nand2_1 _26138_ (.A(\count_instr[5] ),
    .B(_19761_),
    .Y(_04205_));
 sky130_fd_sc_hd__o221a_1 _26139_ (.A1(_18995_),
    .A2(_04130_),
    .B1(_04204_),
    .B2(_19180_),
    .C1(_04205_),
    .X(_01781_));
 sky130_fd_sc_hd__a22o_1 _26140_ (.A1(\irq_mask[5] ),
    .A2(_19739_),
    .B1(_19725_),
    .B2(\timer[5] ),
    .X(_04206_));
 sky130_fd_sc_hd__a21oi_1 _26141_ (.A1(\cpuregs_rs1[5] ),
    .A2(_04190_),
    .B1(_04206_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor2_2 _26142_ (.A(\reg_pc[5] ),
    .B(\decoded_imm[5] ),
    .Y(_04207_));
 sky130_fd_sc_hd__nor2_2 _26143_ (.A(_18859_),
    .B(_20449_),
    .Y(_04208_));
 sky130_fd_sc_hd__nor2_4 _26144_ (.A(_04207_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__o21ai_1 _26145_ (.A1(_04194_),
    .A2(_04199_),
    .B1(_04193_),
    .Y(_04210_));
 sky130_fd_sc_hd__or2_1 _26146_ (.A(_04209_),
    .B(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__nand2_1 _26147_ (.A(_04210_),
    .B(_04209_),
    .Y(_04212_));
 sky130_fd_sc_hd__clkbuf_2 _26148_ (.A(_19090_),
    .X(_04213_));
 sky130_fd_sc_hd__nor2_1 _26149_ (.A(_01784_),
    .B(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__a2bb2o_1 _26150_ (.A1_N(_01778_),
    .A2_N(_20183_),
    .B1(_04162_),
    .B2(_01779_),
    .X(_04215_));
 sky130_fd_sc_hd__a311o_1 _26151_ (.A1(_04211_),
    .A2(_04158_),
    .A3(_04212_),
    .B1(_04214_),
    .C1(_04215_),
    .X(_01785_));
 sky130_vsdinv _26152_ (.A(net61),
    .Y(_01786_));
 sky130_fd_sc_hd__a22o_1 _26153_ (.A1(_04117_),
    .A2(net38),
    .B1(net47),
    .B2(_04119_),
    .X(_04216_));
 sky130_fd_sc_hd__a21oi_1 _26154_ (.A1(net513),
    .A2(_04121_),
    .B1(_04216_),
    .Y(_01787_));
 sky130_fd_sc_hd__o2bb2a_1 _26155_ (.A1_N(_04188_),
    .A2_N(_01789_),
    .B1(_01788_),
    .B2(_20358_),
    .X(_01790_));
 sky130_fd_sc_hd__clkbuf_2 _26156_ (.A(instr_rdinstrh),
    .X(_04217_));
 sky130_fd_sc_hd__nand2_1 _26157_ (.A(\count_instr[38] ),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__o221a_1 _26158_ (.A1(_19053_),
    .A2(_04175_),
    .B1(_04204_),
    .B2(_19212_),
    .C1(_04218_),
    .X(_01794_));
 sky130_fd_sc_hd__nand2_1 _26159_ (.A(\cpuregs_rs1[6] ),
    .B(_04152_),
    .Y(_04219_));
 sky130_fd_sc_hd__o221a_1 _26160_ (.A1(_18382_),
    .A2(_04149_),
    .B1(_04150_),
    .B2(_20373_),
    .C1(_04219_),
    .X(_01796_));
 sky130_fd_sc_hd__nand3_4 _26161_ (.A(_04197_),
    .B(_04195_),
    .C(_04209_),
    .Y(_04220_));
 sky130_fd_sc_hd__o21ba_1 _26162_ (.A1(_04193_),
    .A2(_04207_),
    .B1_N(_04208_),
    .X(_04221_));
 sky130_fd_sc_hd__nand2_1 _26163_ (.A(_20506_),
    .B(_20450_),
    .Y(_04222_));
 sky130_fd_sc_hd__nand2_1 _26164_ (.A(\reg_pc[6] ),
    .B(\decoded_imm[6] ),
    .Y(_04223_));
 sky130_fd_sc_hd__nand2_1 _26165_ (.A(_04222_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__and3_1 _26166_ (.A(_04220_),
    .B(_04221_),
    .C(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__and2_1 _26167_ (.A(_04220_),
    .B(_04221_),
    .X(_04226_));
 sky130_fd_sc_hd__nor2_1 _26168_ (.A(_04224_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__nand2_1 _26169_ (.A(_04141_),
    .B(_01792_),
    .Y(_04228_));
 sky130_fd_sc_hd__o221a_1 _26170_ (.A1(_01791_),
    .A2(_04144_),
    .B1(_19131_),
    .B2(_01797_),
    .C1(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__o31ai_2 _26171_ (.A1(_20194_),
    .A2(_04225_),
    .A3(_04227_),
    .B1(_04229_),
    .Y(_01798_));
 sky130_vsdinv _26172_ (.A(net62),
    .Y(_01799_));
 sky130_fd_sc_hd__a22o_1 _26173_ (.A1(_04117_),
    .A2(net516),
    .B1(net48),
    .B2(_04119_),
    .X(_04230_));
 sky130_fd_sc_hd__a21oi_1 _26174_ (.A1(net57),
    .A2(_04121_),
    .B1(_04230_),
    .Y(_01800_));
 sky130_fd_sc_hd__o2bb2a_1 _26175_ (.A1_N(_04188_),
    .A2_N(_01802_),
    .B1(_01801_),
    .B2(_20358_),
    .X(_01803_));
 sky130_fd_sc_hd__nand2_1 _26176_ (.A(\count_instr[39] ),
    .B(_04217_),
    .Y(_04231_));
 sky130_fd_sc_hd__o221a_1 _26177_ (.A1(_19052_),
    .A2(_04175_),
    .B1(_04204_),
    .B2(_19213_),
    .C1(_04231_),
    .X(_01807_));
 sky130_fd_sc_hd__a22o_1 _26178_ (.A1(\irq_mask[7] ),
    .A2(_19739_),
    .B1(_19725_),
    .B2(\timer[7] ),
    .X(_04232_));
 sky130_fd_sc_hd__a21oi_1 _26179_ (.A1(\cpuregs_rs1[7] ),
    .A2(_04190_),
    .B1(_04232_),
    .Y(_01809_));
 sky130_fd_sc_hd__nor2_1 _26180_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .Y(_04233_));
 sky130_fd_sc_hd__nand2_1 _26181_ (.A(\reg_pc[7] ),
    .B(\decoded_imm[7] ),
    .Y(_04234_));
 sky130_fd_sc_hd__or2b_1 _26182_ (.A(_04233_),
    .B_N(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__o21a_1 _26183_ (.A1(_04224_),
    .A2(_04226_),
    .B1(_04223_),
    .X(_04236_));
 sky130_fd_sc_hd__or2_1 _26184_ (.A(_04235_),
    .B(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_1 _26185_ (.A(_04236_),
    .B(_04235_),
    .Y(_04238_));
 sky130_vsdinv _26186_ (.A(_01804_),
    .Y(_04239_));
 sky130_fd_sc_hd__nor2_1 _26187_ (.A(_01810_),
    .B(_19090_),
    .Y(_04240_));
 sky130_fd_sc_hd__a221o_1 _26188_ (.A1(_18334_),
    .A2(_04239_),
    .B1(_04141_),
    .B2(_01805_),
    .C1(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__a31o_1 _26189_ (.A1(_04237_),
    .A2(_04138_),
    .A3(_04238_),
    .B1(_04241_),
    .X(_01811_));
 sky130_vsdinv _26190_ (.A(net63),
    .Y(_01812_));
 sky130_fd_sc_hd__clkbuf_2 _26191_ (.A(_04112_),
    .X(_04242_));
 sky130_fd_sc_hd__nand2_1 _26192_ (.A(_04242_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_8 _26193_ (.A(latched_is_lb),
    .B(latched_is_lh),
    .Y(_01816_));
 sky130_vsdinv _26194_ (.A(latched_is_lh),
    .Y(_04243_));
 sky130_fd_sc_hd__clkbuf_2 _26195_ (.A(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__nand2_1 _26196_ (.A(_04239_),
    .B(latched_is_lb),
    .Y(_04245_));
 sky130_fd_sc_hd__clkbuf_2 _26197_ (.A(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__o21a_1 _26198_ (.A1(_04244_),
    .A2(_01815_),
    .B1(_04246_),
    .X(_01817_));
 sky130_fd_sc_hd__nand2_1 _26199_ (.A(\count_instr[8] ),
    .B(_19761_),
    .Y(_04247_));
 sky130_fd_sc_hd__o221a_1 _26200_ (.A1(_18915_),
    .A2(_04130_),
    .B1(_04204_),
    .B2(_19287_),
    .C1(_04247_),
    .X(_01821_));
 sky130_fd_sc_hd__nand2_1 _26201_ (.A(\cpuregs_rs1[8] ),
    .B(_04152_),
    .Y(_04248_));
 sky130_fd_sc_hd__o221a_1 _26202_ (.A1(_18406_),
    .A2(_04149_),
    .B1(_04150_),
    .B2(_20412_),
    .C1(_04248_),
    .X(_01823_));
 sky130_fd_sc_hd__nand2_1 _26203_ (.A(_20516_),
    .B(_20452_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_1 _26204_ (.A(\reg_pc[8] ),
    .B(\decoded_imm[8] ),
    .Y(_04250_));
 sky130_fd_sc_hd__nand2_1 _26205_ (.A(_04249_),
    .B(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__o21a_1 _26206_ (.A1(_04223_),
    .A2(_04233_),
    .B1(_04234_),
    .X(_04252_));
 sky130_vsdinv _26207_ (.A(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__or2_1 _26208_ (.A(_04224_),
    .B(_04235_),
    .X(_04254_));
 sky130_fd_sc_hd__a21oi_4 _26209_ (.A1(_04220_),
    .A2(_04221_),
    .B1(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__nor2_1 _26210_ (.A(_04253_),
    .B(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__or2_1 _26211_ (.A(_04251_),
    .B(_04256_),
    .X(_04257_));
 sky130_fd_sc_hd__nand2_1 _26212_ (.A(_04256_),
    .B(_04251_),
    .Y(_04258_));
 sky130_fd_sc_hd__nor2_2 _26213_ (.A(_01818_),
    .B(_20348_),
    .Y(_04259_));
 sky130_fd_sc_hd__a2bb2o_1 _26214_ (.A1_N(_01824_),
    .A2_N(_04142_),
    .B1(_04162_),
    .B2(_01819_),
    .X(_04260_));
 sky130_fd_sc_hd__a311o_1 _26215_ (.A1(_04257_),
    .A2(_04158_),
    .A3(_04258_),
    .B1(_04259_),
    .C1(_04260_),
    .X(_01825_));
 sky130_vsdinv _26216_ (.A(net64),
    .Y(_01826_));
 sky130_fd_sc_hd__nand2_1 _26217_ (.A(_04242_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__o21a_1 _26218_ (.A1(_04244_),
    .A2(_01829_),
    .B1(_04246_),
    .X(_01830_));
 sky130_fd_sc_hd__buf_2 _26219_ (.A(_19760_),
    .X(_04261_));
 sky130_fd_sc_hd__a22o_1 _26220_ (.A1(\count_instr[41] ),
    .A2(_04217_),
    .B1(\count_instr[9] ),
    .B2(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__a21oi_2 _26221_ (.A1(_19763_),
    .A2(\count_cycle[41] ),
    .B1(_04262_),
    .Y(_01834_));
 sky130_fd_sc_hd__a22o_1 _26222_ (.A1(\irq_mask[9] ),
    .A2(_19739_),
    .B1(_19725_),
    .B2(\timer[9] ),
    .X(_04263_));
 sky130_fd_sc_hd__a21oi_1 _26223_ (.A1(\cpuregs_rs1[9] ),
    .A2(_04190_),
    .B1(_04263_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_1 _26224_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .Y(_04264_));
 sky130_fd_sc_hd__nand2_1 _26225_ (.A(\reg_pc[9] ),
    .B(\decoded_imm[9] ),
    .Y(_04265_));
 sky130_fd_sc_hd__or2b_1 _26226_ (.A(_04264_),
    .B_N(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__and2_1 _26227_ (.A(_04257_),
    .B(_04250_),
    .X(_04267_));
 sky130_fd_sc_hd__or2_1 _26228_ (.A(_04266_),
    .B(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__nand2_1 _26229_ (.A(_04267_),
    .B(_04266_),
    .Y(_04269_));
 sky130_fd_sc_hd__nor2_1 _26230_ (.A(_01837_),
    .B(_04213_),
    .Y(_04270_));
 sky130_fd_sc_hd__a2bb2o_1 _26231_ (.A1_N(_01831_),
    .A2_N(_20183_),
    .B1(_04162_),
    .B2(_01832_),
    .X(_04271_));
 sky130_fd_sc_hd__a311o_1 _26232_ (.A1(_04268_),
    .A2(_04158_),
    .A3(_04269_),
    .B1(_04270_),
    .C1(_04271_),
    .X(_01838_));
 sky130_vsdinv _26233_ (.A(net34),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _26234_ (.A(_04242_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o21a_1 _26235_ (.A1(_04244_),
    .A2(_01842_),
    .B1(_04246_),
    .X(_01843_));
 sky130_fd_sc_hd__nand2_1 _26236_ (.A(\count_instr[42] ),
    .B(_04217_),
    .Y(_04272_));
 sky130_fd_sc_hd__o221a_1 _26237_ (.A1(_19050_),
    .A2(_04175_),
    .B1(_04204_),
    .B2(_19277_),
    .C1(_04272_),
    .X(_01847_));
 sky130_vsdinv _26238_ (.A(\timer[10] ),
    .Y(_04273_));
 sky130_fd_sc_hd__clkbuf_2 _26239_ (.A(_04151_),
    .X(_04274_));
 sky130_fd_sc_hd__nand2_1 _26240_ (.A(\cpuregs_rs1[10] ),
    .B(_04274_),
    .Y(_04275_));
 sky130_fd_sc_hd__o221a_1 _26241_ (.A1(_18405_),
    .A2(_04149_),
    .B1(_04150_),
    .B2(_04273_),
    .C1(_04275_),
    .X(_01849_));
 sky130_fd_sc_hd__nor2_2 _26242_ (.A(\reg_pc[10] ),
    .B(\decoded_imm[10] ),
    .Y(_04276_));
 sky130_fd_sc_hd__nor2_4 _26243_ (.A(_20530_),
    .B(_20455_),
    .Y(_04277_));
 sky130_fd_sc_hd__or2_1 _26244_ (.A(_04276_),
    .B(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__or2_1 _26245_ (.A(_04251_),
    .B(_04266_),
    .X(_04279_));
 sky130_fd_sc_hd__o21bai_4 _26246_ (.A1(_04253_),
    .A2(_04255_),
    .B1_N(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__o21a_1 _26247_ (.A1(_04250_),
    .A2(_04264_),
    .B1(_04265_),
    .X(_04281_));
 sky130_fd_sc_hd__and2_1 _26248_ (.A(_04280_),
    .B(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__or2_1 _26249_ (.A(_04278_),
    .B(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__nand2_1 _26250_ (.A(_04282_),
    .B(_04278_),
    .Y(_04284_));
 sky130_fd_sc_hd__o22ai_4 _26251_ (.A1(_01844_),
    .A2(_04144_),
    .B1(_04142_),
    .B2(_01850_),
    .Y(_04285_));
 sky130_fd_sc_hd__a21o_1 _26252_ (.A1(_04122_),
    .A2(_01845_),
    .B1(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__a31o_1 _26253_ (.A1(_04283_),
    .A2(_04138_),
    .A3(_04284_),
    .B1(_04286_),
    .X(_01851_));
 sky130_vsdinv _26254_ (.A(net35),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _26255_ (.A(_04242_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__o21a_1 _26256_ (.A1(_04244_),
    .A2(_01855_),
    .B1(_04246_),
    .X(_01856_));
 sky130_fd_sc_hd__nand2_1 _26257_ (.A(\count_instr[11] ),
    .B(_19761_),
    .Y(_04287_));
 sky130_fd_sc_hd__o221a_1 _26258_ (.A1(_18981_),
    .A2(_04130_),
    .B1(_04204_),
    .B2(_19281_),
    .C1(_04287_),
    .X(_01860_));
 sky130_fd_sc_hd__clkbuf_2 _26259_ (.A(_18494_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_2 _26260_ (.A(_18492_),
    .X(_04289_));
 sky130_fd_sc_hd__nand2_1 _26261_ (.A(\cpuregs_rs1[11] ),
    .B(_04274_),
    .Y(_04290_));
 sky130_fd_sc_hd__o221a_2 _26262_ (.A1(_18408_),
    .A2(_04288_),
    .B1(_04289_),
    .B2(_20379_),
    .C1(_04290_),
    .X(_01862_));
 sky130_fd_sc_hd__nor2_2 _26263_ (.A(_20540_),
    .B(_20456_),
    .Y(_04291_));
 sky130_fd_sc_hd__nor2_1 _26264_ (.A(\reg_pc[11] ),
    .B(\decoded_imm[11] ),
    .Y(_04292_));
 sky130_fd_sc_hd__a21oi_4 _26265_ (.A1(_04280_),
    .A2(_04281_),
    .B1(_04276_),
    .Y(_04293_));
 sky130_fd_sc_hd__nor2_1 _26266_ (.A(_04277_),
    .B(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__or3_2 _26267_ (.A(_04291_),
    .B(_04292_),
    .C(_04294_),
    .X(_04295_));
 sky130_fd_sc_hd__o21ai_1 _26268_ (.A1(_04291_),
    .A2(_04292_),
    .B1(_04294_),
    .Y(_04296_));
 sky130_fd_sc_hd__buf_2 _26269_ (.A(_20150_),
    .X(_04297_));
 sky130_fd_sc_hd__o22a_1 _26270_ (.A1(_01857_),
    .A2(_20182_),
    .B1(_19106_),
    .B2(_01863_),
    .X(_04298_));
 sky130_fd_sc_hd__a21bo_1 _26271_ (.A1(_04297_),
    .A2(_01858_),
    .B1_N(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__a31o_1 _26272_ (.A1(_04295_),
    .A2(_04138_),
    .A3(_04296_),
    .B1(_04299_),
    .X(_01864_));
 sky130_vsdinv _26273_ (.A(net517),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _26274_ (.A(_04242_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__o21a_1 _26275_ (.A1(_04244_),
    .A2(_01868_),
    .B1(_04246_),
    .X(_01869_));
 sky130_fd_sc_hd__nand2_1 _26276_ (.A(_19763_),
    .B(\count_cycle[44] ),
    .Y(_04300_));
 sky130_fd_sc_hd__o221a_1 _26277_ (.A1(_18876_),
    .A2(_04130_),
    .B1(_19066_),
    .B2(_04132_),
    .C1(_04300_),
    .X(_01873_));
 sky130_fd_sc_hd__clkbuf_2 _26278_ (.A(_18493_),
    .X(_04301_));
 sky130_fd_sc_hd__a22o_1 _26279_ (.A1(\irq_mask[12] ),
    .A2(_04301_),
    .B1(_19725_),
    .B2(\timer[12] ),
    .X(_04302_));
 sky130_fd_sc_hd__a21oi_2 _26280_ (.A1(\cpuregs_rs1[12] ),
    .A2(_04190_),
    .B1(_04302_),
    .Y(_01875_));
 sky130_fd_sc_hd__clkbuf_4 _26281_ (.A(_19090_),
    .X(_04303_));
 sky130_fd_sc_hd__o22ai_4 _26282_ (.A1(_01870_),
    .A2(_20348_),
    .B1(_04303_),
    .B2(_01876_),
    .Y(_04304_));
 sky130_fd_sc_hd__nor2_1 _26283_ (.A(\reg_pc[12] ),
    .B(\decoded_imm[12] ),
    .Y(_04305_));
 sky130_fd_sc_hd__nor2_4 _26284_ (.A(_20548_),
    .B(_20457_),
    .Y(_04306_));
 sky130_fd_sc_hd__or2_1 _26285_ (.A(_04305_),
    .B(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__o22ai_4 _26286_ (.A1(\reg_pc[11] ),
    .A2(\decoded_imm[11] ),
    .B1(_04277_),
    .B2(_04293_),
    .Y(_04308_));
 sky130_vsdinv _26287_ (.A(_04291_),
    .Y(_04309_));
 sky130_fd_sc_hd__nand2_1 _26288_ (.A(_04308_),
    .B(_04309_),
    .Y(_04310_));
 sky130_vsdinv _26289_ (.A(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__or2_1 _26290_ (.A(_04307_),
    .B(_04311_),
    .X(_04312_));
 sky130_fd_sc_hd__nand2_1 _26291_ (.A(_04311_),
    .B(_04307_),
    .Y(_04313_));
 sky130_fd_sc_hd__and3_1 _26292_ (.A(_04312_),
    .B(\cpu_state[4] ),
    .C(_04313_),
    .X(_04314_));
 sky130_fd_sc_hd__a211o_1 _26293_ (.A1(_04122_),
    .A2(_01871_),
    .B1(_04304_),
    .C1(_04314_),
    .X(_01877_));
 sky130_vsdinv _26294_ (.A(net37),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _26295_ (.A(_04242_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__o21a_1 _26296_ (.A1(_04244_),
    .A2(_01881_),
    .B1(_04246_),
    .X(_01882_));
 sky130_fd_sc_hd__buf_2 _26297_ (.A(_04129_),
    .X(_04315_));
 sky130_fd_sc_hd__buf_2 _26298_ (.A(_04133_),
    .X(_04316_));
 sky130_fd_sc_hd__nand2_1 _26299_ (.A(\count_instr[13] ),
    .B(_19761_),
    .Y(_04317_));
 sky130_fd_sc_hd__o221a_1 _26300_ (.A1(_18875_),
    .A2(_04315_),
    .B1(_04316_),
    .B2(_19218_),
    .C1(_04317_),
    .X(_01886_));
 sky130_fd_sc_hd__clkbuf_2 _26301_ (.A(instr_timer),
    .X(_04318_));
 sky130_fd_sc_hd__a22o_1 _26302_ (.A1(\irq_mask[13] ),
    .A2(_04301_),
    .B1(_04318_),
    .B2(\timer[13] ),
    .X(_04319_));
 sky130_fd_sc_hd__a21oi_4 _26303_ (.A1(\cpuregs_rs1[13] ),
    .A2(_04190_),
    .B1(_04319_),
    .Y(_01888_));
 sky130_fd_sc_hd__nor2_2 _26304_ (.A(_20555_),
    .B(_20458_),
    .Y(_04320_));
 sky130_fd_sc_hd__nor2_1 _26305_ (.A(\reg_pc[13] ),
    .B(\decoded_imm[13] ),
    .Y(_04321_));
 sky130_fd_sc_hd__a22oi_4 _26306_ (.A1(_20548_),
    .A2(_20457_),
    .B1(_04308_),
    .B2(_04309_),
    .Y(_04322_));
 sky130_fd_sc_hd__nor2_1 _26307_ (.A(_04306_),
    .B(_04322_),
    .Y(_04323_));
 sky130_fd_sc_hd__or3_1 _26308_ (.A(_04320_),
    .B(_04321_),
    .C(_04323_),
    .X(_04324_));
 sky130_fd_sc_hd__o21ai_1 _26309_ (.A1(_04320_),
    .A2(_04321_),
    .B1(_04323_),
    .Y(_04325_));
 sky130_fd_sc_hd__o22a_1 _26310_ (.A1(_01883_),
    .A2(_20182_),
    .B1(_19106_),
    .B2(_01889_),
    .X(_04326_));
 sky130_fd_sc_hd__a21bo_1 _26311_ (.A1(_04297_),
    .A2(_01884_),
    .B1_N(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__a31o_1 _26312_ (.A1(_04324_),
    .A2(_04138_),
    .A3(_04325_),
    .B1(_04327_),
    .X(_01890_));
 sky130_vsdinv _26313_ (.A(net38),
    .Y(_01891_));
 sky130_fd_sc_hd__nand2_1 _26314_ (.A(_04128_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hd__o21a_1 _26315_ (.A1(_04243_),
    .A2(_01894_),
    .B1(_04245_),
    .X(_01895_));
 sky130_fd_sc_hd__nand2_1 _26316_ (.A(\count_instr[14] ),
    .B(_04261_),
    .Y(_04328_));
 sky130_fd_sc_hd__o221a_1 _26317_ (.A1(_18968_),
    .A2(_04315_),
    .B1(_04316_),
    .B2(_19219_),
    .C1(_04328_),
    .X(_01899_));
 sky130_fd_sc_hd__nand2_1 _26318_ (.A(\cpuregs_rs1[14] ),
    .B(_04274_),
    .Y(_04329_));
 sky130_fd_sc_hd__o221a_1 _26319_ (.A1(_18428_),
    .A2(_04288_),
    .B1(_04289_),
    .B2(_20383_),
    .C1(_04329_),
    .X(_01901_));
 sky130_fd_sc_hd__clkbuf_4 _26320_ (.A(_20182_),
    .X(_04330_));
 sky130_fd_sc_hd__o22ai_4 _26321_ (.A1(_01896_),
    .A2(_04330_),
    .B1(_04303_),
    .B2(_01902_),
    .Y(_04331_));
 sky130_fd_sc_hd__nor2_1 _26322_ (.A(\reg_pc[14] ),
    .B(\decoded_imm[14] ),
    .Y(_04332_));
 sky130_fd_sc_hd__nor2_4 _26323_ (.A(_20562_),
    .B(_20459_),
    .Y(_04333_));
 sky130_fd_sc_hd__or2_1 _26324_ (.A(_04332_),
    .B(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__o22ai_4 _26325_ (.A1(\reg_pc[13] ),
    .A2(\decoded_imm[13] ),
    .B1(_04306_),
    .B2(_04322_),
    .Y(_04335_));
 sky130_vsdinv _26326_ (.A(_04320_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _26327_ (.A(_04335_),
    .B(_04336_),
    .Y(_04337_));
 sky130_vsdinv _26328_ (.A(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__or2_1 _26329_ (.A(_04334_),
    .B(_04338_),
    .X(_04339_));
 sky130_fd_sc_hd__nand2_1 _26330_ (.A(_04338_),
    .B(_04334_),
    .Y(_04340_));
 sky130_fd_sc_hd__and3_1 _26331_ (.A(_04339_),
    .B(\cpu_state[4] ),
    .C(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__a211o_1 _26332_ (.A1(_04122_),
    .A2(_01897_),
    .B1(_04331_),
    .C1(_04341_),
    .X(_01903_));
 sky130_vsdinv _26333_ (.A(net516),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_1 _26334_ (.A(_04128_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__o21a_4 _26335_ (.A1(_04243_),
    .A2(_01907_),
    .B1(_04245_),
    .X(_01908_));
 sky130_fd_sc_hd__nand2_1 _26336_ (.A(\count_instr[15] ),
    .B(_04261_),
    .Y(_04342_));
 sky130_fd_sc_hd__o221a_1 _26337_ (.A1(_18967_),
    .A2(_04315_),
    .B1(_04316_),
    .B2(_19220_),
    .C1(_04342_),
    .X(_01912_));
 sky130_fd_sc_hd__nand2_1 _26338_ (.A(\cpuregs_rs1[15] ),
    .B(_04274_),
    .Y(_04343_));
 sky130_fd_sc_hd__o221a_1 _26339_ (.A1(_18603_),
    .A2(_04288_),
    .B1(_04289_),
    .B2(_20382_),
    .C1(_04343_),
    .X(_01914_));
 sky130_fd_sc_hd__nor2_2 _26340_ (.A(_20568_),
    .B(_20460_),
    .Y(_04344_));
 sky130_vsdinv _26341_ (.A(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__nand2_1 _26342_ (.A(_20568_),
    .B(_20460_),
    .Y(_04346_));
 sky130_fd_sc_hd__nand2_1 _26343_ (.A(_04345_),
    .B(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__a22oi_4 _26344_ (.A1(_20562_),
    .A2(_20459_),
    .B1(_04335_),
    .B2(_04336_),
    .Y(_04348_));
 sky130_fd_sc_hd__nor2_2 _26345_ (.A(_04333_),
    .B(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__nor2_2 _26346_ (.A(_04347_),
    .B(_04349_),
    .Y(_04350_));
 sky130_fd_sc_hd__nor2_1 _26347_ (.A(_20194_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__nand2_1 _26348_ (.A(_04349_),
    .B(_04347_),
    .Y(_04352_));
 sky130_fd_sc_hd__o22ai_4 _26349_ (.A1(_01909_),
    .A2(_04330_),
    .B1(_19091_),
    .B2(_01915_),
    .Y(_04353_));
 sky130_fd_sc_hd__a221o_1 _26350_ (.A1(_04122_),
    .A2(_01910_),
    .B1(_04351_),
    .B2(_04352_),
    .C1(_04353_),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_1 _26351_ (.A(net431),
    .B(net40),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _26352_ (.A(_19763_),
    .B(\count_cycle[48] ),
    .Y(_04354_));
 sky130_fd_sc_hd__o221a_1 _26353_ (.A1(_18874_),
    .A2(_04315_),
    .B1(_19044_),
    .B2(_04132_),
    .C1(_04354_),
    .X(_01921_));
 sky130_fd_sc_hd__buf_2 _26354_ (.A(_04151_),
    .X(_04355_));
 sky130_fd_sc_hd__a22o_1 _26355_ (.A1(\irq_mask[16] ),
    .A2(_04301_),
    .B1(_04318_),
    .B2(\timer[16] ),
    .X(_04356_));
 sky130_fd_sc_hd__a21oi_4 _26356_ (.A1(\cpuregs_rs1[16] ),
    .A2(_04355_),
    .B1(_04356_),
    .Y(_01923_));
 sky130_fd_sc_hd__o22ai_4 _26357_ (.A1(\reg_pc[15] ),
    .A2(\decoded_imm[15] ),
    .B1(_04333_),
    .B2(_04348_),
    .Y(_04357_));
 sky130_fd_sc_hd__nor2_2 _26358_ (.A(_20575_),
    .B(_20462_),
    .Y(_04358_));
 sky130_vsdinv _26359_ (.A(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__nand2_1 _26360_ (.A(_20575_),
    .B(_20462_),
    .Y(_04360_));
 sky130_fd_sc_hd__nand2_2 _26361_ (.A(_04359_),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__and3_1 _26362_ (.A(_04357_),
    .B(_04345_),
    .C(_04361_),
    .X(_04362_));
 sky130_fd_sc_hd__nor2_2 _26363_ (.A(_04344_),
    .B(_04350_),
    .Y(_04363_));
 sky130_fd_sc_hd__nor2_4 _26364_ (.A(_04361_),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__nand2_1 _26365_ (.A(_04162_),
    .B(_01919_),
    .Y(_04365_));
 sky130_fd_sc_hd__o221a_2 _26366_ (.A1(_01918_),
    .A2(_04144_),
    .B1(_04142_),
    .B2(_01924_),
    .C1(_04365_),
    .X(_04366_));
 sky130_fd_sc_hd__o31ai_4 _26367_ (.A1(_20194_),
    .A2(_04362_),
    .A3(_04364_),
    .B1(_04366_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2_1 _26368_ (.A(net431),
    .B(net41),
    .Y(_01926_));
 sky130_fd_sc_hd__nand2_1 _26369_ (.A(\count_instr[49] ),
    .B(_04217_),
    .Y(_04367_));
 sky130_fd_sc_hd__o221a_1 _26370_ (.A1(_19036_),
    .A2(_04175_),
    .B1(_04316_),
    .B2(_19224_),
    .C1(_04367_),
    .X(_01930_));
 sky130_fd_sc_hd__a22o_1 _26371_ (.A1(\irq_mask[17] ),
    .A2(_04301_),
    .B1(_04318_),
    .B2(\timer[17] ),
    .X(_04368_));
 sky130_fd_sc_hd__a21oi_1 _26372_ (.A1(\cpuregs_rs1[17] ),
    .A2(_04355_),
    .B1(_04368_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_2 _26373_ (.A(\reg_pc[17] ),
    .B(\decoded_imm[17] ),
    .Y(_04369_));
 sky130_fd_sc_hd__nor2_1 _26374_ (.A(_20580_),
    .B(_20463_),
    .Y(_04370_));
 sky130_fd_sc_hd__nor2_1 _26375_ (.A(_04369_),
    .B(_04370_),
    .Y(_04371_));
 sky130_vsdinv _26376_ (.A(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__nor2_1 _26377_ (.A(_04358_),
    .B(_04364_),
    .Y(_04373_));
 sky130_fd_sc_hd__or2_1 _26378_ (.A(_04372_),
    .B(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__nand2_1 _26379_ (.A(_04373_),
    .B(_04372_),
    .Y(_04375_));
 sky130_fd_sc_hd__nor2_2 _26380_ (.A(_01933_),
    .B(_04213_),
    .Y(_04376_));
 sky130_fd_sc_hd__clkbuf_2 _26381_ (.A(_20150_),
    .X(_04377_));
 sky130_fd_sc_hd__a2bb2o_2 _26382_ (.A1_N(_01927_),
    .A2_N(_20183_),
    .B1(_04377_),
    .B2(_01928_),
    .X(_04378_));
 sky130_fd_sc_hd__a311o_1 _26383_ (.A1(_04374_),
    .A2(_04158_),
    .A3(_04375_),
    .B1(_04376_),
    .C1(_04378_),
    .X(_01934_));
 sky130_fd_sc_hd__nand2_1 _26384_ (.A(net431),
    .B(net42),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2_1 _26385_ (.A(\count_instr[18] ),
    .B(_04261_),
    .Y(_04379_));
 sky130_fd_sc_hd__o221a_1 _26386_ (.A1(_18964_),
    .A2(_04315_),
    .B1(_04316_),
    .B2(_19225_),
    .C1(_04379_),
    .X(_01939_));
 sky130_vsdinv _26387_ (.A(\timer[18] ),
    .Y(_04380_));
 sky130_fd_sc_hd__nand2_1 _26388_ (.A(\cpuregs_rs1[18] ),
    .B(_04274_),
    .Y(_04381_));
 sky130_fd_sc_hd__o221a_1 _26389_ (.A1(_18394_),
    .A2(_04288_),
    .B1(_04289_),
    .B2(_04380_),
    .C1(_04381_),
    .X(_01941_));
 sky130_fd_sc_hd__nand2_1 _26390_ (.A(_20586_),
    .B(_20464_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_2 _26391_ (.A(\reg_pc[18] ),
    .B(\decoded_imm[18] ),
    .Y(_04383_));
 sky130_fd_sc_hd__nand2_1 _26392_ (.A(_04382_),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__o21bai_4 _26393_ (.A1(_04369_),
    .A2(_04359_),
    .B1_N(_04370_),
    .Y(_04385_));
 sky130_fd_sc_hd__or2_1 _26394_ (.A(_04361_),
    .B(_04372_),
    .X(_04386_));
 sky130_fd_sc_hd__a21oi_4 _26395_ (.A1(_04357_),
    .A2(_04345_),
    .B1(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__nor2_1 _26396_ (.A(_04385_),
    .B(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__or2_1 _26397_ (.A(_04384_),
    .B(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__nand2_1 _26398_ (.A(_04388_),
    .B(_04384_),
    .Y(_04390_));
 sky130_fd_sc_hd__o22a_1 _26399_ (.A1(_01936_),
    .A2(_18328_),
    .B1(_19106_),
    .B2(_01942_),
    .X(_04391_));
 sky130_fd_sc_hd__a21bo_1 _26400_ (.A1(_04297_),
    .A2(_01937_),
    .B1_N(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__a31o_1 _26401_ (.A1(_04389_),
    .A2(_04171_),
    .A3(_04390_),
    .B1(_04392_),
    .X(_01943_));
 sky130_fd_sc_hd__nand2_1 _26402_ (.A(net431),
    .B(net515),
    .Y(_01944_));
 sky130_vsdinv _26403_ (.A(\count_cycle[19] ),
    .Y(_01947_));
 sky130_fd_sc_hd__clkbuf_2 _26404_ (.A(instr_rdcycleh),
    .X(_04393_));
 sky130_fd_sc_hd__nand2_1 _26405_ (.A(_04393_),
    .B(\count_cycle[51] ),
    .Y(_04394_));
 sky130_fd_sc_hd__o221a_1 _26406_ (.A1(_18921_),
    .A2(_04315_),
    .B1(_18901_),
    .B2(_04132_),
    .C1(_04394_),
    .X(_01948_));
 sky130_fd_sc_hd__a22o_1 _26407_ (.A1(\irq_mask[19] ),
    .A2(_04301_),
    .B1(_04318_),
    .B2(\timer[19] ),
    .X(_04395_));
 sky130_fd_sc_hd__a21oi_1 _26408_ (.A1(\cpuregs_rs1[19] ),
    .A2(_04355_),
    .B1(_04395_),
    .Y(_01950_));
 sky130_fd_sc_hd__nor2_2 _26409_ (.A(_20595_),
    .B(_20465_),
    .Y(_04396_));
 sky130_vsdinv _26410_ (.A(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _26411_ (.A(_20595_),
    .B(_20465_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand2_1 _26412_ (.A(_04397_),
    .B(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__o22ai_4 _26413_ (.A1(\reg_pc[18] ),
    .A2(\decoded_imm[18] ),
    .B1(_04385_),
    .B2(_04387_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand2_1 _26414_ (.A(_04400_),
    .B(_04383_),
    .Y(_04401_));
 sky130_vsdinv _26415_ (.A(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__or2_1 _26416_ (.A(_04399_),
    .B(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__nand2_1 _26417_ (.A(_04402_),
    .B(_04399_),
    .Y(_04404_));
 sky130_fd_sc_hd__nor2_1 _26418_ (.A(_01951_),
    .B(_04213_),
    .Y(_04405_));
 sky130_fd_sc_hd__buf_1 _26419_ (.A(_20182_),
    .X(_04406_));
 sky130_fd_sc_hd__a2bb2o_2 _26420_ (.A1_N(_01945_),
    .A2_N(_04406_),
    .B1(_04377_),
    .B2(_01946_),
    .X(_04407_));
 sky130_fd_sc_hd__a311o_1 _26421_ (.A1(_04403_),
    .A2(_04158_),
    .A3(_04404_),
    .B1(_04405_),
    .C1(_04407_),
    .X(_01952_));
 sky130_fd_sc_hd__nand2_1 _26422_ (.A(net432),
    .B(net514),
    .Y(_01953_));
 sky130_fd_sc_hd__clkbuf_2 _26423_ (.A(_04129_),
    .X(_04408_));
 sky130_fd_sc_hd__nand2_1 _26424_ (.A(\count_instr[20] ),
    .B(_04261_),
    .Y(_04409_));
 sky130_fd_sc_hd__o221a_1 _26425_ (.A1(_18920_),
    .A2(_04408_),
    .B1(_04316_),
    .B2(_19257_),
    .C1(_04409_),
    .X(_01957_));
 sky130_fd_sc_hd__nand2_1 _26426_ (.A(\cpuregs_rs1[20] ),
    .B(_04274_),
    .Y(_04410_));
 sky130_fd_sc_hd__o221a_1 _26427_ (.A1(_18425_),
    .A2(_04288_),
    .B1(_04289_),
    .B2(_20390_),
    .C1(_04410_),
    .X(_01959_));
 sky130_vsdinv _26428_ (.A(_01955_),
    .Y(_04411_));
 sky130_fd_sc_hd__a22oi_4 _26429_ (.A1(_20595_),
    .A2(_20465_),
    .B1(_04400_),
    .B2(_04383_),
    .Y(_04412_));
 sky130_vsdinv _26430_ (.A(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__nor2_1 _26431_ (.A(\reg_pc[20] ),
    .B(\decoded_imm[20] ),
    .Y(_04414_));
 sky130_fd_sc_hd__nor2_2 _26432_ (.A(_20601_),
    .B(_20466_),
    .Y(_04415_));
 sky130_fd_sc_hd__or2_2 _26433_ (.A(_04414_),
    .B(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__and3_1 _26434_ (.A(_04413_),
    .B(_04397_),
    .C(_04416_),
    .X(_04417_));
 sky130_fd_sc_hd__a21oi_4 _26435_ (.A1(_04413_),
    .A2(_04397_),
    .B1(_04416_),
    .Y(_04418_));
 sky130_fd_sc_hd__o32a_2 _26436_ (.A1(_18487_),
    .A2(_04417_),
    .A3(_04418_),
    .B1(_04330_),
    .B2(_01954_),
    .X(_04419_));
 sky130_fd_sc_hd__o221ai_4 _26437_ (.A1(_04160_),
    .A2(_01960_),
    .B1(_18520_),
    .B2(_04411_),
    .C1(_04419_),
    .Y(_01961_));
 sky130_fd_sc_hd__clkbuf_2 _26438_ (.A(_04114_),
    .X(_04420_));
 sky130_fd_sc_hd__nand2_1 _26439_ (.A(_04420_),
    .B(net46),
    .Y(_01962_));
 sky130_fd_sc_hd__a22o_1 _26440_ (.A1(\count_instr[53] ),
    .A2(instr_rdinstrh),
    .B1(\count_instr[21] ),
    .B2(_19760_),
    .X(_04421_));
 sky130_fd_sc_hd__a21oi_2 _26441_ (.A1(_19763_),
    .A2(\count_cycle[53] ),
    .B1(_04421_),
    .Y(_01966_));
 sky130_vsdinv _26442_ (.A(\timer[21] ),
    .Y(_04422_));
 sky130_fd_sc_hd__clkbuf_2 _26443_ (.A(_04151_),
    .X(_04423_));
 sky130_fd_sc_hd__nand2_1 _26444_ (.A(\cpuregs_rs1[21] ),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__o221a_1 _26445_ (.A1(_18421_),
    .A2(_04288_),
    .B1(_04289_),
    .B2(_04422_),
    .C1(_04424_),
    .X(_01968_));
 sky130_fd_sc_hd__nor2_1 _26446_ (.A(\reg_pc[21] ),
    .B(\decoded_imm[21] ),
    .Y(_04425_));
 sky130_fd_sc_hd__nor2_4 _26447_ (.A(_20609_),
    .B(_20467_),
    .Y(_04426_));
 sky130_fd_sc_hd__nor2_1 _26448_ (.A(_04425_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__or3_1 _26449_ (.A(_04415_),
    .B(_04427_),
    .C(_04418_),
    .X(_04428_));
 sky130_fd_sc_hd__o21ai_1 _26450_ (.A1(_04415_),
    .A2(_04418_),
    .B1(_04427_),
    .Y(_04429_));
 sky130_fd_sc_hd__nor2_1 _26451_ (.A(_01969_),
    .B(_04213_),
    .Y(_04430_));
 sky130_fd_sc_hd__a2bb2o_1 _26452_ (.A1_N(_01963_),
    .A2_N(_04406_),
    .B1(_04377_),
    .B2(_01964_),
    .X(_04431_));
 sky130_fd_sc_hd__a311o_1 _26453_ (.A1(_04428_),
    .A2(_18479_),
    .A3(_04429_),
    .B1(_04430_),
    .C1(_04431_),
    .X(_01970_));
 sky130_fd_sc_hd__nand2_1 _26454_ (.A(_04420_),
    .B(net47),
    .Y(_01971_));
 sky130_fd_sc_hd__nand2_1 _26455_ (.A(_04393_),
    .B(\count_cycle[54] ),
    .Y(_04432_));
 sky130_fd_sc_hd__o221a_1 _26456_ (.A1(_18950_),
    .A2(_04408_),
    .B1(_18905_),
    .B2(_04132_),
    .C1(_04432_),
    .X(_01975_));
 sky130_fd_sc_hd__a22o_1 _26457_ (.A1(\irq_mask[22] ),
    .A2(_04301_),
    .B1(_04318_),
    .B2(\timer[22] ),
    .X(_04433_));
 sky130_fd_sc_hd__a21oi_1 _26458_ (.A1(\cpuregs_rs1[22] ),
    .A2(_04355_),
    .B1(_04433_),
    .Y(_01977_));
 sky130_fd_sc_hd__o22ai_4 _26459_ (.A1(\reg_pc[20] ),
    .A2(\decoded_imm[20] ),
    .B1(_04396_),
    .B2(_04412_),
    .Y(_04434_));
 sky130_vsdinv _26460_ (.A(_04415_),
    .Y(_04435_));
 sky130_fd_sc_hd__a22oi_4 _26461_ (.A1(_20609_),
    .A2(_20467_),
    .B1(_04434_),
    .B2(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hd__nor2_1 _26462_ (.A(\reg_pc[22] ),
    .B(\decoded_imm[22] ),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_2 _26463_ (.A(_20614_),
    .B(_20469_),
    .Y(_04438_));
 sky130_fd_sc_hd__or2_1 _26464_ (.A(_04437_),
    .B(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__or3b_2 _26465_ (.A(_04426_),
    .B(_04436_),
    .C_N(_04439_),
    .X(_04440_));
 sky130_vsdinv _26466_ (.A(_04436_),
    .Y(_04441_));
 sky130_vsdinv _26467_ (.A(_04426_),
    .Y(_04442_));
 sky130_fd_sc_hd__a21o_1 _26468_ (.A1(_04441_),
    .A2(_04442_),
    .B1(_04439_),
    .X(_04443_));
 sky130_fd_sc_hd__nor2_1 _26469_ (.A(_01978_),
    .B(_04213_),
    .Y(_04444_));
 sky130_fd_sc_hd__a2bb2o_1 _26470_ (.A1_N(_01972_),
    .A2_N(_04406_),
    .B1(_04377_),
    .B2(_01973_),
    .X(_04445_));
 sky130_fd_sc_hd__a311o_2 _26471_ (.A1(_04440_),
    .A2(_04443_),
    .A3(_04171_),
    .B1(_04444_),
    .C1(_04445_),
    .X(_01979_));
 sky130_fd_sc_hd__nand2_1 _26472_ (.A(_04420_),
    .B(net48),
    .Y(_01980_));
 sky130_fd_sc_hd__nand2_1 _26473_ (.A(_04393_),
    .B(\count_cycle[55] ),
    .Y(_04446_));
 sky130_fd_sc_hd__o221a_1 _26474_ (.A1(_18954_),
    .A2(_04408_),
    .B1(_18904_),
    .B2(_04132_),
    .C1(_04446_),
    .X(_01984_));
 sky130_fd_sc_hd__a22o_1 _26475_ (.A1(\irq_mask[23] ),
    .A2(_18493_),
    .B1(_04318_),
    .B2(\timer[23] ),
    .X(_04447_));
 sky130_fd_sc_hd__a21oi_1 _26476_ (.A1(\cpuregs_rs1[23] ),
    .A2(_04355_),
    .B1(_04447_),
    .Y(_01986_));
 sky130_fd_sc_hd__nor2_1 _26477_ (.A(\reg_pc[23] ),
    .B(\decoded_imm[23] ),
    .Y(_04448_));
 sky130_fd_sc_hd__nor2_2 _26478_ (.A(_20622_),
    .B(_20470_),
    .Y(_04449_));
 sky130_fd_sc_hd__nor2_1 _26479_ (.A(_04448_),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__o22ai_4 _26480_ (.A1(\reg_pc[22] ),
    .A2(\decoded_imm[22] ),
    .B1(_04426_),
    .B2(_04436_),
    .Y(_04451_));
 sky130_vsdinv _26481_ (.A(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__or3_1 _26482_ (.A(_04438_),
    .B(_04450_),
    .C(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__o21ai_1 _26483_ (.A1(_04438_),
    .A2(_04452_),
    .B1(_04450_),
    .Y(_04454_));
 sky130_fd_sc_hd__nor2_1 _26484_ (.A(_01987_),
    .B(_04303_),
    .Y(_04455_));
 sky130_fd_sc_hd__a2bb2o_1 _26485_ (.A1_N(_01981_),
    .A2_N(_04406_),
    .B1(_04377_),
    .B2(_01982_),
    .X(_04456_));
 sky130_fd_sc_hd__a311o_2 _26486_ (.A1(_04453_),
    .A2(_18479_),
    .A3(_04454_),
    .B1(_04455_),
    .C1(_04456_),
    .X(_01988_));
 sky130_fd_sc_hd__nand2_1 _26487_ (.A(_04420_),
    .B(net49),
    .Y(_01989_));
 sky130_fd_sc_hd__nand2_1 _26488_ (.A(_04393_),
    .B(\count_cycle[56] ),
    .Y(_04457_));
 sky130_fd_sc_hd__o221a_1 _26489_ (.A1(_18944_),
    .A2(_04408_),
    .B1(_19024_),
    .B2(_04135_),
    .C1(_04457_),
    .X(_01993_));
 sky130_fd_sc_hd__clkbuf_2 _26490_ (.A(_18494_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_2 _26491_ (.A(_18492_),
    .X(_04459_));
 sky130_fd_sc_hd__nand2_1 _26492_ (.A(\cpuregs_rs1[24] ),
    .B(_04423_),
    .Y(_04460_));
 sky130_fd_sc_hd__o221a_1 _26493_ (.A1(_18398_),
    .A2(_04458_),
    .B1(_04459_),
    .B2(_20435_),
    .C1(_04460_),
    .X(_01995_));
 sky130_fd_sc_hd__o2bb2a_1 _26494_ (.A1_N(_04297_),
    .A2_N(_01991_),
    .B1(_01996_),
    .B2(_04142_),
    .X(_04461_));
 sky130_vsdinv _26495_ (.A(_04449_),
    .Y(_04462_));
 sky130_fd_sc_hd__nor2_1 _26496_ (.A(_20628_),
    .B(_20471_),
    .Y(_04463_));
 sky130_vsdinv _26497_ (.A(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_1 _26498_ (.A(_20628_),
    .B(_20471_),
    .Y(_04465_));
 sky130_fd_sc_hd__nand2_1 _26499_ (.A(_04464_),
    .B(_04465_),
    .Y(_04466_));
 sky130_vsdinv _26500_ (.A(_04438_),
    .Y(_04467_));
 sky130_fd_sc_hd__a22oi_4 _26501_ (.A1(_20622_),
    .A2(_20470_),
    .B1(_04451_),
    .B2(_04467_),
    .Y(_04468_));
 sky130_vsdinv _26502_ (.A(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hd__a21o_1 _26503_ (.A1(_04469_),
    .A2(_04462_),
    .B1(_04466_),
    .X(_04470_));
 sky130_vsdinv _26504_ (.A(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__a311o_2 _26505_ (.A1(_04462_),
    .A2(_04454_),
    .A3(_04466_),
    .B1(_20194_),
    .C1(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__o211ai_4 _26506_ (.A1(_20348_),
    .A2(_01990_),
    .B1(_04461_),
    .C1(_04472_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand2_1 _26507_ (.A(_04420_),
    .B(net50),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_1 _26508_ (.A(\count_instr[57] ),
    .B(_04217_),
    .Y(_04473_));
 sky130_fd_sc_hd__o221a_1 _26509_ (.A1(_18884_),
    .A2(_04131_),
    .B1(_04133_),
    .B2(_19244_),
    .C1(_04473_),
    .X(_02002_));
 sky130_fd_sc_hd__a22o_1 _26510_ (.A1(\irq_mask[25] ),
    .A2(_18493_),
    .B1(instr_timer),
    .B2(\timer[25] ),
    .X(_04474_));
 sky130_fd_sc_hd__a21oi_1 _26511_ (.A1(\cpuregs_rs1[25] ),
    .A2(_04355_),
    .B1(_04474_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_1 _26512_ (.A(\reg_pc[25] ),
    .B(\decoded_imm[25] ),
    .Y(_04475_));
 sky130_fd_sc_hd__nor2_1 _26513_ (.A(_20637_),
    .B(_20472_),
    .Y(_04476_));
 sky130_fd_sc_hd__nor2_1 _26514_ (.A(_04475_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__or3_1 _26515_ (.A(_04463_),
    .B(_04477_),
    .C(_04471_),
    .X(_04478_));
 sky130_vsdinv _26516_ (.A(_04477_),
    .Y(_04479_));
 sky130_fd_sc_hd__a21o_1 _26517_ (.A1(_04470_),
    .A2(_04464_),
    .B1(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__nor2_1 _26518_ (.A(_02005_),
    .B(_04303_),
    .Y(_04481_));
 sky130_fd_sc_hd__a2bb2o_1 _26519_ (.A1_N(_01999_),
    .A2_N(_04406_),
    .B1(_04377_),
    .B2(_02000_),
    .X(_04482_));
 sky130_fd_sc_hd__a311o_2 _26520_ (.A1(_04478_),
    .A2(_18479_),
    .A3(_04480_),
    .B1(_04481_),
    .C1(_04482_),
    .X(_02006_));
 sky130_fd_sc_hd__nand2_1 _26521_ (.A(_04420_),
    .B(net51),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2_1 _26522_ (.A(_04393_),
    .B(\count_cycle[58] ),
    .Y(_04483_));
 sky130_fd_sc_hd__o221a_1 _26523_ (.A1(_18871_),
    .A2(_04408_),
    .B1(_18883_),
    .B2(_04135_),
    .C1(_04483_),
    .X(_02011_));
 sky130_vsdinv _26524_ (.A(\timer[26] ),
    .Y(_04484_));
 sky130_fd_sc_hd__nand2_1 _26525_ (.A(\cpuregs_rs1[26] ),
    .B(_04423_),
    .Y(_04485_));
 sky130_fd_sc_hd__o221a_1 _26526_ (.A1(_18400_),
    .A2(_04458_),
    .B1(_04459_),
    .B2(_04484_),
    .C1(_04485_),
    .X(_02013_));
 sky130_fd_sc_hd__or2_1 _26527_ (.A(_04466_),
    .B(_04479_),
    .X(_04486_));
 sky130_fd_sc_hd__o21bai_2 _26528_ (.A1(_04449_),
    .A2(_04468_),
    .B1_N(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__o21ba_1 _26529_ (.A1(_04475_),
    .A2(_04464_),
    .B1_N(_04476_),
    .X(_04488_));
 sky130_fd_sc_hd__nand2_1 _26530_ (.A(_20643_),
    .B(_20473_),
    .Y(_04489_));
 sky130_fd_sc_hd__nand2_1 _26531_ (.A(\reg_pc[26] ),
    .B(\decoded_imm[26] ),
    .Y(_04490_));
 sky130_fd_sc_hd__nand2_1 _26532_ (.A(_04489_),
    .B(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__a21o_1 _26533_ (.A1(_04487_),
    .A2(_04488_),
    .B1(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__nand3_1 _26534_ (.A(_04487_),
    .B(_04488_),
    .C(_04491_),
    .Y(_04493_));
 sky130_fd_sc_hd__o22ai_1 _26535_ (.A1(_02008_),
    .A2(_04144_),
    .B1(_04142_),
    .B2(_02014_),
    .Y(_04494_));
 sky130_fd_sc_hd__a21o_1 _26536_ (.A1(_04297_),
    .A2(_02009_),
    .B1(_04494_),
    .X(_04495_));
 sky130_fd_sc_hd__a31o_1 _26537_ (.A1(_04492_),
    .A2(_04171_),
    .A3(_04493_),
    .B1(_04495_),
    .X(_02015_));
 sky130_fd_sc_hd__clkbuf_4 _26538_ (.A(_04114_),
    .X(_04496_));
 sky130_fd_sc_hd__nand2_1 _26539_ (.A(_04496_),
    .B(net52),
    .Y(_02016_));
 sky130_vsdinv _26540_ (.A(\count_cycle[27] ),
    .Y(_02019_));
 sky130_fd_sc_hd__a22o_1 _26541_ (.A1(_18927_),
    .A2(instr_rdinstrh),
    .B1(\count_instr[27] ),
    .B2(_19760_),
    .X(_04497_));
 sky130_fd_sc_hd__a21oi_1 _26542_ (.A1(_19763_),
    .A2(\count_cycle[59] ),
    .B1(_04497_),
    .Y(_02020_));
 sky130_vsdinv _26543_ (.A(\timer[27] ),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_1 _26544_ (.A(\cpuregs_rs1[27] ),
    .B(_04423_),
    .Y(_04499_));
 sky130_fd_sc_hd__o221a_1 _26545_ (.A1(_18402_),
    .A2(_04458_),
    .B1(_04459_),
    .B2(_04498_),
    .C1(_04499_),
    .X(_02022_));
 sky130_fd_sc_hd__nor2_2 _26546_ (.A(\reg_pc[27] ),
    .B(\decoded_imm[27] ),
    .Y(_04500_));
 sky130_fd_sc_hd__nor2_2 _26547_ (.A(_20653_),
    .B(_20474_),
    .Y(_04501_));
 sky130_fd_sc_hd__nor2_1 _26548_ (.A(_04500_),
    .B(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand2_1 _26549_ (.A(_04492_),
    .B(_04490_),
    .Y(_04503_));
 sky130_fd_sc_hd__or2_1 _26550_ (.A(_04502_),
    .B(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__nand2_1 _26551_ (.A(_04503_),
    .B(_04502_),
    .Y(_04505_));
 sky130_fd_sc_hd__o22a_1 _26552_ (.A1(_02017_),
    .A2(_18328_),
    .B1(_19106_),
    .B2(_02023_),
    .X(_04506_));
 sky130_fd_sc_hd__a21bo_1 _26553_ (.A1(_04297_),
    .A2(_02018_),
    .B1_N(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__a31o_1 _26554_ (.A1(_04504_),
    .A2(_04171_),
    .A3(_04505_),
    .B1(_04507_),
    .X(_02024_));
 sky130_fd_sc_hd__nand2_1 _26555_ (.A(_04496_),
    .B(net53),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_1 _26556_ (.A(_04393_),
    .B(\count_cycle[60] ),
    .Y(_04508_));
 sky130_fd_sc_hd__o221a_1 _26557_ (.A1(_18939_),
    .A2(_04408_),
    .B1(_19008_),
    .B2(_04135_),
    .C1(_04508_),
    .X(_02029_));
 sky130_fd_sc_hd__nand2_1 _26558_ (.A(\cpuregs_rs1[28] ),
    .B(_04423_),
    .Y(_04509_));
 sky130_fd_sc_hd__o221a_1 _26559_ (.A1(_18435_),
    .A2(_04458_),
    .B1(_04459_),
    .B2(_20443_),
    .C1(_04509_),
    .X(_02031_));
 sky130_fd_sc_hd__o21ba_1 _26560_ (.A1(_04490_),
    .A2(_04500_),
    .B1_N(_04501_),
    .X(_04510_));
 sky130_vsdinv _26561_ (.A(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__or3_4 _26562_ (.A(_04500_),
    .B(_04501_),
    .C(_04491_),
    .X(_04512_));
 sky130_fd_sc_hd__a21oi_4 _26563_ (.A1(_04487_),
    .A2(_04488_),
    .B1(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__nor2_1 _26564_ (.A(_20659_),
    .B(_20475_),
    .Y(_04514_));
 sky130_vsdinv _26565_ (.A(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__nand2_1 _26566_ (.A(_20659_),
    .B(_20475_),
    .Y(_04516_));
 sky130_fd_sc_hd__nand2_1 _26567_ (.A(_04515_),
    .B(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__or3b_2 _26568_ (.A(_04511_),
    .B(_04513_),
    .C_N(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__o21bai_1 _26569_ (.A1(_04511_),
    .A2(_04513_),
    .B1_N(_04517_),
    .Y(_04519_));
 sky130_fd_sc_hd__nor2_1 _26570_ (.A(_02032_),
    .B(_04303_),
    .Y(_04520_));
 sky130_fd_sc_hd__a2bb2o_1 _26571_ (.A1_N(_02026_),
    .A2_N(_04406_),
    .B1(_20150_),
    .B2(_02027_),
    .X(_04521_));
 sky130_fd_sc_hd__a311o_1 _26572_ (.A1(_04518_),
    .A2(_18479_),
    .A3(_04519_),
    .B1(_04520_),
    .C1(_04521_),
    .X(_02033_));
 sky130_fd_sc_hd__nand2_1 _26573_ (.A(_04496_),
    .B(net54),
    .Y(_02034_));
 sky130_fd_sc_hd__a22o_1 _26574_ (.A1(\count_instr[29] ),
    .A2(_19760_),
    .B1(instr_rdcycleh),
    .B2(\count_cycle[61] ),
    .X(_04522_));
 sky130_fd_sc_hd__a21oi_1 _26575_ (.A1(\count_instr[61] ),
    .A2(_19752_),
    .B1(_04522_),
    .Y(_02038_));
 sky130_fd_sc_hd__a22o_1 _26576_ (.A1(\irq_mask[29] ),
    .A2(_18493_),
    .B1(instr_timer),
    .B2(\timer[29] ),
    .X(_04523_));
 sky130_fd_sc_hd__a21oi_1 _26577_ (.A1(\cpuregs_rs1[29] ),
    .A2(_04152_),
    .B1(_04523_),
    .Y(_02040_));
 sky130_vsdinv _26578_ (.A(_02036_),
    .Y(_04524_));
 sky130_fd_sc_hd__o22ai_4 _26579_ (.A1(\reg_pc[28] ),
    .A2(\decoded_imm[28] ),
    .B1(_04511_),
    .B2(_04513_),
    .Y(_04525_));
 sky130_fd_sc_hd__nor2_1 _26580_ (.A(\reg_pc[29] ),
    .B(\decoded_imm[29] ),
    .Y(_04526_));
 sky130_fd_sc_hd__nor2_1 _26581_ (.A(_20669_),
    .B(_20476_),
    .Y(_04527_));
 sky130_fd_sc_hd__or2_1 _26582_ (.A(_04526_),
    .B(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__a21oi_1 _26583_ (.A1(_04525_),
    .A2(_04515_),
    .B1(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__and3_1 _26584_ (.A(_04525_),
    .B(_04515_),
    .C(_04528_),
    .X(_04530_));
 sky130_fd_sc_hd__o32a_2 _26585_ (.A1(_18487_),
    .A2(_04529_),
    .A3(_04530_),
    .B1(_04330_),
    .B2(_02035_),
    .X(_04531_));
 sky130_fd_sc_hd__o221ai_4 _26586_ (.A1(_04160_),
    .A2(_02041_),
    .B1(_18520_),
    .B2(_04524_),
    .C1(_04531_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_1 _26587_ (.A(_04496_),
    .B(net513),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _26588_ (.A(instr_rdcycleh),
    .B(\count_cycle[62] ),
    .Y(_04532_));
 sky130_fd_sc_hd__o221a_1 _26589_ (.A1(_18931_),
    .A2(_04129_),
    .B1(_19013_),
    .B2(_04135_),
    .C1(_04532_),
    .X(_02047_));
 sky130_fd_sc_hd__nand2_1 _26590_ (.A(\cpuregs_rs1[30] ),
    .B(_04423_),
    .Y(_04533_));
 sky130_fd_sc_hd__o221a_1 _26591_ (.A1(_18434_),
    .A2(_04458_),
    .B1(_04459_),
    .B2(_20401_),
    .C1(_04533_),
    .X(_02049_));
 sky130_fd_sc_hd__nand2_2 _26592_ (.A(\reg_pc[30] ),
    .B(\decoded_imm[30] ),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_2 _26593_ (.A(_20676_),
    .B(_20477_),
    .Y(_04535_));
 sky130_fd_sc_hd__a22oi_2 _26594_ (.A1(_20669_),
    .A2(_20476_),
    .B1(_04525_),
    .B2(_04515_),
    .Y(_04536_));
 sky130_fd_sc_hd__a211o_1 _26595_ (.A1(_04534_),
    .A2(_04535_),
    .B1(_04527_),
    .C1(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__nand2_1 _26596_ (.A(_04535_),
    .B(_04534_),
    .Y(_04538_));
 sky130_fd_sc_hd__o21bai_1 _26597_ (.A1(_04527_),
    .A2(_04536_),
    .B1_N(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__nand2_1 _26598_ (.A(_04141_),
    .B(_02045_),
    .Y(_04540_));
 sky130_fd_sc_hd__o221ai_2 _26599_ (.A1(_02044_),
    .A2(_04330_),
    .B1(_02050_),
    .B2(_04303_),
    .C1(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a31o_1 _26600_ (.A1(_04537_),
    .A2(_04171_),
    .A3(_04539_),
    .B1(_04541_),
    .X(_02051_));
 sky130_fd_sc_hd__nand2_1 _26601_ (.A(_04496_),
    .B(net57),
    .Y(_02052_));
 sky130_fd_sc_hd__nand2_1 _26602_ (.A(\count_instr[31] ),
    .B(_04261_),
    .Y(_04542_));
 sky130_fd_sc_hd__o221a_1 _26603_ (.A1(_18930_),
    .A2(_04129_),
    .B1(_04133_),
    .B2(_19175_),
    .C1(_04542_),
    .X(_02056_));
 sky130_fd_sc_hd__nand2_1 _26604_ (.A(\cpuregs_rs1[31] ),
    .B(_04151_),
    .Y(_04543_));
 sky130_fd_sc_hd__o221a_1 _26605_ (.A1(_18438_),
    .A2(_04458_),
    .B1(_04459_),
    .B2(_20400_),
    .C1(_04543_),
    .X(_02058_));
 sky130_fd_sc_hd__xnor2_1 _26606_ (.A(\reg_pc[31] ),
    .B(\decoded_imm[31] ),
    .Y(_04544_));
 sky130_fd_sc_hd__a21oi_1 _26607_ (.A1(_04539_),
    .A2(_04534_),
    .B1(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand3_1 _26608_ (.A(_04539_),
    .B(_04534_),
    .C(_04544_),
    .Y(_04546_));
 sky130_fd_sc_hd__nand2_1 _26609_ (.A(_04546_),
    .B(_18479_),
    .Y(_04547_));
 sky130_fd_sc_hd__nand2_1 _26610_ (.A(_04141_),
    .B(_02054_),
    .Y(_04548_));
 sky130_fd_sc_hd__o221ai_1 _26611_ (.A1(_02053_),
    .A2(_04330_),
    .B1(_02059_),
    .B2(_19091_),
    .C1(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__o21bai_2 _26612_ (.A1(_04545_),
    .A2(_04547_),
    .B1_N(_04549_),
    .Y(_02060_));
 sky130_fd_sc_hd__or2_1 _26613_ (.A(\decoded_rd[4] ),
    .B(_00308_),
    .X(_02061_));
 sky130_fd_sc_hd__o21ai_1 _26614_ (.A1(_02064_),
    .A2(_20195_),
    .B1(_04160_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor3_1 _26615_ (.A(_19162_),
    .B(_02410_),
    .C(_00308_),
    .Y(_02066_));
 sky130_fd_sc_hd__and3_1 _26616_ (.A(_18498_),
    .B(_20194_),
    .C(_20348_),
    .X(_02067_));
 sky130_fd_sc_hd__nand2_1 _26617_ (.A(is_beq_bne_blt_bge_bltu_bgeu),
    .B(_00343_),
    .Y(_04550_));
 sky130_fd_sc_hd__a211o_1 _26618_ (.A1(_04550_),
    .A2(_04138_),
    .B1(_18496_),
    .C1(_18334_),
    .X(_02068_));
 sky130_fd_sc_hd__and2_2 _26619_ (.A(_18343_),
    .B(latched_store),
    .X(_04551_));
 sky130_fd_sc_hd__buf_4 _26620_ (.A(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__nor2_8 _26621_ (.A(_18536_),
    .B(_04552_),
    .Y(_02069_));
 sky130_fd_sc_hd__nor2_1 _26622_ (.A(_20355_),
    .B(_20480_),
    .Y(_04553_));
 sky130_fd_sc_hd__a221o_1 _26623_ (.A1(_18415_),
    .A2(_18530_),
    .B1(_04552_),
    .B2(_02070_),
    .C1(_04553_),
    .X(_02071_));
 sky130_fd_sc_hd__buf_2 _26624_ (.A(_18530_),
    .X(_04554_));
 sky130_fd_sc_hd__and3_1 _26625_ (.A(_18344_),
    .B(_18486_),
    .C(_01465_),
    .X(_04555_));
 sky130_fd_sc_hd__a221o_1 _26626_ (.A1(_20692_),
    .A2(\reg_next_pc[1] ),
    .B1(_04554_),
    .B2(_18417_),
    .C1(_04555_),
    .X(_02072_));
 sky130_fd_sc_hd__buf_1 _26627_ (.A(_18529_),
    .X(_04556_));
 sky130_fd_sc_hd__and3_1 _26628_ (.A(_18623_),
    .B(_04556_),
    .C(\irq_pending[2] ),
    .X(_04557_));
 sky130_fd_sc_hd__a221o_1 _26629_ (.A1(_20692_),
    .A2(\reg_next_pc[2] ),
    .B1(_04552_),
    .B2(_00293_),
    .C1(_04557_),
    .X(_02074_));
 sky130_fd_sc_hd__nand2_1 _26630_ (.A(_20489_),
    .B(_02073_),
    .Y(_04558_));
 sky130_fd_sc_hd__nand2_1 _26631_ (.A(\reg_pc[3] ),
    .B(\reg_pc[2] ),
    .Y(_04559_));
 sky130_fd_sc_hd__and2_1 _26632_ (.A(_04558_),
    .B(_04559_),
    .X(_02075_));
 sky130_fd_sc_hd__and3_1 _26633_ (.A(_18418_),
    .B(_04556_),
    .C(\irq_pending[3] ),
    .X(_04560_));
 sky130_fd_sc_hd__a221o_1 _26634_ (.A1(_20692_),
    .A2(\reg_next_pc[3] ),
    .B1(_04552_),
    .B2(_01468_),
    .C1(_04560_),
    .X(_02076_));
 sky130_fd_sc_hd__or2_1 _26635_ (.A(_04559_),
    .B(_20495_),
    .X(_04561_));
 sky130_fd_sc_hd__nand2_1 _26636_ (.A(_20495_),
    .B(_04559_),
    .Y(_04562_));
 sky130_fd_sc_hd__and2_1 _26637_ (.A(_04561_),
    .B(_04562_),
    .X(_02077_));
 sky130_fd_sc_hd__nor2_1 _26638_ (.A(_20355_),
    .B(_01471_),
    .Y(_04563_));
 sky130_fd_sc_hd__a221o_1 _26639_ (.A1(_18384_),
    .A2(_18530_),
    .B1(_04552_),
    .B2(_01472_),
    .C1(_04563_),
    .X(_02078_));
 sky130_fd_sc_hd__nor2_2 _26640_ (.A(_18859_),
    .B(_04561_),
    .Y(_04564_));
 sky130_fd_sc_hd__and2_1 _26641_ (.A(_04561_),
    .B(_18859_),
    .X(_04565_));
 sky130_fd_sc_hd__nor2_1 _26642_ (.A(_04564_),
    .B(_04565_),
    .Y(_02079_));
 sky130_fd_sc_hd__and3_1 _26643_ (.A(_18385_),
    .B(_04556_),
    .C(\irq_pending[5] ),
    .X(_04566_));
 sky130_fd_sc_hd__a221o_1 _26644_ (.A1(_20692_),
    .A2(\reg_next_pc[5] ),
    .B1(_04552_),
    .B2(_01476_),
    .C1(_04566_),
    .X(_02080_));
 sky130_fd_sc_hd__nor2_1 _26645_ (.A(\reg_pc[6] ),
    .B(_04564_),
    .Y(_04567_));
 sky130_fd_sc_hd__and2_1 _26646_ (.A(_04564_),
    .B(\reg_pc[6] ),
    .X(_04568_));
 sky130_fd_sc_hd__nor2_1 _26647_ (.A(_04567_),
    .B(_04568_),
    .Y(_02081_));
 sky130_fd_sc_hd__buf_2 _26648_ (.A(_04551_),
    .X(_04569_));
 sky130_fd_sc_hd__and3_1 _26649_ (.A(_18382_),
    .B(_04556_),
    .C(\irq_pending[6] ),
    .X(_04570_));
 sky130_fd_sc_hd__a221o_1 _26650_ (.A1(_20692_),
    .A2(\reg_next_pc[6] ),
    .B1(_04569_),
    .B2(_01479_),
    .C1(_04570_),
    .X(_02082_));
 sky130_fd_sc_hd__or2_1 _26651_ (.A(\reg_pc[7] ),
    .B(_04568_),
    .X(_04571_));
 sky130_fd_sc_hd__nand2_2 _26652_ (.A(_04568_),
    .B(\reg_pc[7] ),
    .Y(_04572_));
 sky130_fd_sc_hd__and2_1 _26653_ (.A(_04571_),
    .B(_04572_),
    .X(_02083_));
 sky130_fd_sc_hd__buf_2 _26654_ (.A(_18526_),
    .X(_04573_));
 sky130_fd_sc_hd__and3_1 _26655_ (.A(_18387_),
    .B(_04556_),
    .C(\irq_pending[7] ),
    .X(_04574_));
 sky130_fd_sc_hd__a221o_1 _26656_ (.A1(_04573_),
    .A2(\reg_next_pc[7] ),
    .B1(_04569_),
    .B2(_01482_),
    .C1(_04574_),
    .X(_02084_));
 sky130_fd_sc_hd__nor2_2 _26657_ (.A(_20516_),
    .B(_04572_),
    .Y(_04575_));
 sky130_fd_sc_hd__and2_1 _26658_ (.A(_04572_),
    .B(_20516_),
    .X(_04576_));
 sky130_fd_sc_hd__nor2_1 _26659_ (.A(_04575_),
    .B(_04576_),
    .Y(_02085_));
 sky130_fd_sc_hd__and3_1 _26660_ (.A(_18406_),
    .B(_04556_),
    .C(\irq_pending[8] ),
    .X(_04577_));
 sky130_fd_sc_hd__a221o_1 _26661_ (.A1(_04573_),
    .A2(\reg_next_pc[8] ),
    .B1(_04569_),
    .B2(_01485_),
    .C1(_04577_),
    .X(_02086_));
 sky130_fd_sc_hd__nor2_1 _26662_ (.A(\reg_pc[9] ),
    .B(_04575_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand2_1 _26663_ (.A(_04575_),
    .B(\reg_pc[9] ),
    .Y(_04579_));
 sky130_vsdinv _26664_ (.A(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__nor2_1 _26665_ (.A(_04578_),
    .B(_04580_),
    .Y(_02087_));
 sky130_fd_sc_hd__buf_2 _26666_ (.A(_18525_),
    .X(_04581_));
 sky130_fd_sc_hd__and3_1 _26667_ (.A(_18344_),
    .B(_18486_),
    .C(_01488_),
    .X(_04582_));
 sky130_fd_sc_hd__a221o_1 _26668_ (.A1(_04554_),
    .A2(_18407_),
    .B1(_04581_),
    .B2(\reg_next_pc[9] ),
    .C1(_04582_),
    .X(_02088_));
 sky130_fd_sc_hd__nor2_2 _26669_ (.A(_20530_),
    .B(_04579_),
    .Y(_04583_));
 sky130_fd_sc_hd__nor2_1 _26670_ (.A(\reg_pc[10] ),
    .B(_04580_),
    .Y(_04584_));
 sky130_fd_sc_hd__nor2_1 _26671_ (.A(_04583_),
    .B(_04584_),
    .Y(_02089_));
 sky130_fd_sc_hd__buf_1 _26672_ (.A(\irq_state[1] ),
    .X(_04585_));
 sky130_fd_sc_hd__and3_1 _26673_ (.A(_18405_),
    .B(_04585_),
    .C(\irq_pending[10] ),
    .X(_04586_));
 sky130_fd_sc_hd__a221o_1 _26674_ (.A1(_04573_),
    .A2(\reg_next_pc[10] ),
    .B1(_04569_),
    .B2(_01491_),
    .C1(_04586_),
    .X(_02090_));
 sky130_fd_sc_hd__or2_1 _26675_ (.A(\reg_pc[11] ),
    .B(_04583_),
    .X(_04587_));
 sky130_fd_sc_hd__nand2_1 _26676_ (.A(_04583_),
    .B(\reg_pc[11] ),
    .Y(_04588_));
 sky130_fd_sc_hd__and2_1 _26677_ (.A(_04587_),
    .B(_04588_),
    .X(_02091_));
 sky130_fd_sc_hd__and3_1 _26678_ (.A(_18408_),
    .B(_04585_),
    .C(\irq_pending[11] ),
    .X(_04589_));
 sky130_fd_sc_hd__a221o_1 _26679_ (.A1(_04573_),
    .A2(\reg_next_pc[11] ),
    .B1(_04569_),
    .B2(_01494_),
    .C1(_04589_),
    .X(_02092_));
 sky130_fd_sc_hd__nor2_1 _26680_ (.A(_20548_),
    .B(_04588_),
    .Y(_04590_));
 sky130_fd_sc_hd__and2_1 _26681_ (.A(_04588_),
    .B(_20548_),
    .X(_04591_));
 sky130_fd_sc_hd__nor2_1 _26682_ (.A(_04590_),
    .B(_04591_),
    .Y(_02093_));
 sky130_fd_sc_hd__and3_1 _26683_ (.A(_18429_),
    .B(_04585_),
    .C(\irq_pending[12] ),
    .X(_04592_));
 sky130_fd_sc_hd__a221o_1 _26684_ (.A1(_04573_),
    .A2(\reg_next_pc[12] ),
    .B1(_04569_),
    .B2(_01497_),
    .C1(_04592_),
    .X(_02094_));
 sky130_fd_sc_hd__nor2_1 _26685_ (.A(\reg_pc[13] ),
    .B(_04590_),
    .Y(_04593_));
 sky130_fd_sc_hd__and2_1 _26686_ (.A(_04590_),
    .B(\reg_pc[13] ),
    .X(_04594_));
 sky130_fd_sc_hd__nor2_1 _26687_ (.A(_04593_),
    .B(_04594_),
    .Y(_02095_));
 sky130_fd_sc_hd__and3_1 _26688_ (.A(_18344_),
    .B(_18486_),
    .C(_01500_),
    .X(_04595_));
 sky130_fd_sc_hd__a221o_1 _26689_ (.A1(_04573_),
    .A2(\reg_next_pc[13] ),
    .B1(_04554_),
    .B2(_18430_),
    .C1(_04595_),
    .X(_02096_));
 sky130_fd_sc_hd__or2_1 _26690_ (.A(\reg_pc[14] ),
    .B(_04594_),
    .X(_04596_));
 sky130_fd_sc_hd__nand2_1 _26691_ (.A(_04594_),
    .B(\reg_pc[14] ),
    .Y(_04597_));
 sky130_fd_sc_hd__and2_1 _26692_ (.A(_04596_),
    .B(_04597_),
    .X(_02097_));
 sky130_fd_sc_hd__clkbuf_2 _26693_ (.A(_18526_),
    .X(_04598_));
 sky130_fd_sc_hd__clkbuf_2 _26694_ (.A(_04551_),
    .X(_04599_));
 sky130_fd_sc_hd__and3_1 _26695_ (.A(_18428_),
    .B(_04585_),
    .C(\irq_pending[14] ),
    .X(_04600_));
 sky130_fd_sc_hd__a221o_1 _26696_ (.A1(_04598_),
    .A2(\reg_next_pc[14] ),
    .B1(_04599_),
    .B2(_01503_),
    .C1(_04600_),
    .X(_02098_));
 sky130_fd_sc_hd__nor2_2 _26697_ (.A(_20568_),
    .B(_04597_),
    .Y(_04601_));
 sky130_fd_sc_hd__and2_1 _26698_ (.A(_04597_),
    .B(_20568_),
    .X(_04602_));
 sky130_fd_sc_hd__nor2_1 _26699_ (.A(_04601_),
    .B(_04602_),
    .Y(_02099_));
 sky130_fd_sc_hd__and3_1 _26700_ (.A(_18344_),
    .B(_18485_),
    .C(_01506_),
    .X(_04603_));
 sky130_fd_sc_hd__a221o_1 _26701_ (.A1(_04554_),
    .A2(_18431_),
    .B1(_04581_),
    .B2(\reg_next_pc[15] ),
    .C1(_04603_),
    .X(_02100_));
 sky130_fd_sc_hd__or2_1 _26702_ (.A(\reg_pc[16] ),
    .B(_04601_),
    .X(_04604_));
 sky130_fd_sc_hd__nand2_2 _26703_ (.A(_04601_),
    .B(\reg_pc[16] ),
    .Y(_04605_));
 sky130_fd_sc_hd__and2_1 _26704_ (.A(_04604_),
    .B(_04605_),
    .X(_02101_));
 sky130_fd_sc_hd__and3_1 _26705_ (.A(_18343_),
    .B(_18485_),
    .C(_01509_),
    .X(_04606_));
 sky130_fd_sc_hd__a221o_1 _26706_ (.A1(_04598_),
    .A2(\reg_next_pc[16] ),
    .B1(_18530_),
    .B2(_18393_),
    .C1(_04606_),
    .X(_02102_));
 sky130_fd_sc_hd__nor2_4 _26707_ (.A(_20580_),
    .B(_04605_),
    .Y(_04607_));
 sky130_fd_sc_hd__and2_1 _26708_ (.A(_04605_),
    .B(_20580_),
    .X(_04608_));
 sky130_fd_sc_hd__nor2_1 _26709_ (.A(_04607_),
    .B(_04608_),
    .Y(_02103_));
 sky130_fd_sc_hd__and3_1 _26710_ (.A(_18390_),
    .B(_04585_),
    .C(\irq_pending[17] ),
    .X(_04609_));
 sky130_fd_sc_hd__a221o_1 _26711_ (.A1(_04598_),
    .A2(\reg_next_pc[17] ),
    .B1(_04599_),
    .B2(_01512_),
    .C1(_04609_),
    .X(_02104_));
 sky130_fd_sc_hd__nor2_1 _26712_ (.A(\reg_pc[18] ),
    .B(_04607_),
    .Y(_04610_));
 sky130_fd_sc_hd__nand2_1 _26713_ (.A(_04607_),
    .B(\reg_pc[18] ),
    .Y(_04611_));
 sky130_vsdinv _26714_ (.A(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_1 _26715_ (.A(_04610_),
    .B(_04612_),
    .Y(_02105_));
 sky130_fd_sc_hd__and3_1 _26716_ (.A(_18394_),
    .B(_04585_),
    .C(\irq_pending[18] ),
    .X(_04613_));
 sky130_fd_sc_hd__a221o_1 _26717_ (.A1(_04598_),
    .A2(\reg_next_pc[18] ),
    .B1(_04599_),
    .B2(_01515_),
    .C1(_04613_),
    .X(_02106_));
 sky130_fd_sc_hd__nor2_1 _26718_ (.A(_20595_),
    .B(_04611_),
    .Y(_04614_));
 sky130_fd_sc_hd__nor2_1 _26719_ (.A(\reg_pc[19] ),
    .B(_04612_),
    .Y(_04615_));
 sky130_fd_sc_hd__nor2_1 _26720_ (.A(_04614_),
    .B(_04615_),
    .Y(_02107_));
 sky130_fd_sc_hd__and3_1 _26721_ (.A(_18343_),
    .B(_18485_),
    .C(_01518_),
    .X(_04616_));
 sky130_fd_sc_hd__a221o_1 _26722_ (.A1(_04554_),
    .A2(_18391_),
    .B1(_04581_),
    .B2(\reg_next_pc[19] ),
    .C1(_04616_),
    .X(_02108_));
 sky130_fd_sc_hd__or2_1 _26723_ (.A(\reg_pc[20] ),
    .B(_04614_),
    .X(_04617_));
 sky130_fd_sc_hd__nand2_1 _26724_ (.A(_04614_),
    .B(\reg_pc[20] ),
    .Y(_04618_));
 sky130_fd_sc_hd__and2_1 _26725_ (.A(_04617_),
    .B(_04618_),
    .X(_02109_));
 sky130_fd_sc_hd__buf_1 _26726_ (.A(\irq_state[1] ),
    .X(_04619_));
 sky130_fd_sc_hd__and3_1 _26727_ (.A(_18425_),
    .B(_04619_),
    .C(\irq_pending[20] ),
    .X(_04620_));
 sky130_fd_sc_hd__a221o_1 _26728_ (.A1(_04598_),
    .A2(\reg_next_pc[20] ),
    .B1(_04599_),
    .B2(_01521_),
    .C1(_04620_),
    .X(_02110_));
 sky130_fd_sc_hd__nor2_2 _26729_ (.A(_20609_),
    .B(_04618_),
    .Y(_04621_));
 sky130_fd_sc_hd__and2_1 _26730_ (.A(_04618_),
    .B(_20609_),
    .X(_04622_));
 sky130_fd_sc_hd__nor2_1 _26731_ (.A(_04621_),
    .B(_04622_),
    .Y(_02111_));
 sky130_fd_sc_hd__and3_1 _26732_ (.A(_18421_),
    .B(_04619_),
    .C(\irq_pending[21] ),
    .X(_04623_));
 sky130_fd_sc_hd__a221o_1 _26733_ (.A1(_04598_),
    .A2(\reg_next_pc[21] ),
    .B1(_04599_),
    .B2(_01524_),
    .C1(_04623_),
    .X(_02112_));
 sky130_fd_sc_hd__nor2_1 _26734_ (.A(\reg_pc[22] ),
    .B(_04621_),
    .Y(_04624_));
 sky130_fd_sc_hd__nand2_1 _26735_ (.A(_04621_),
    .B(\reg_pc[22] ),
    .Y(_04625_));
 sky130_vsdinv _26736_ (.A(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__nor2_1 _26737_ (.A(_04624_),
    .B(_04626_),
    .Y(_02113_));
 sky130_fd_sc_hd__and3_1 _26738_ (.A(_18343_),
    .B(_18485_),
    .C(_01527_),
    .X(_04627_));
 sky130_fd_sc_hd__a221o_1 _26739_ (.A1(_04554_),
    .A2(_18422_),
    .B1(_18526_),
    .B2(\reg_next_pc[22] ),
    .C1(_04627_),
    .X(_02114_));
 sky130_fd_sc_hd__nor2_2 _26740_ (.A(_20622_),
    .B(_04625_),
    .Y(_04628_));
 sky130_fd_sc_hd__nor2_1 _26741_ (.A(\reg_pc[23] ),
    .B(_04626_),
    .Y(_04629_));
 sky130_fd_sc_hd__nor2_1 _26742_ (.A(_04628_),
    .B(_04629_),
    .Y(_02115_));
 sky130_fd_sc_hd__buf_2 _26743_ (.A(_18525_),
    .X(_04630_));
 sky130_fd_sc_hd__and3_1 _26744_ (.A(_18423_),
    .B(_04619_),
    .C(\irq_pending[23] ),
    .X(_04631_));
 sky130_fd_sc_hd__a221o_1 _26745_ (.A1(_04630_),
    .A2(\reg_next_pc[23] ),
    .B1(_04599_),
    .B2(_01530_),
    .C1(_04631_),
    .X(_02116_));
 sky130_fd_sc_hd__or2_1 _26746_ (.A(\reg_pc[24] ),
    .B(_04628_),
    .X(_04632_));
 sky130_fd_sc_hd__nand2_1 _26747_ (.A(_04628_),
    .B(\reg_pc[24] ),
    .Y(_04633_));
 sky130_fd_sc_hd__and2_1 _26748_ (.A(_04632_),
    .B(_04633_),
    .X(_02117_));
 sky130_fd_sc_hd__buf_2 _26749_ (.A(_04551_),
    .X(_04634_));
 sky130_fd_sc_hd__and3_1 _26750_ (.A(_18398_),
    .B(_04619_),
    .C(\irq_pending[24] ),
    .X(_04635_));
 sky130_fd_sc_hd__a221o_1 _26751_ (.A1(_04630_),
    .A2(\reg_next_pc[24] ),
    .B1(_04634_),
    .B2(_01533_),
    .C1(_04635_),
    .X(_02118_));
 sky130_fd_sc_hd__or2_2 _26752_ (.A(_20637_),
    .B(_04633_),
    .X(_04636_));
 sky130_fd_sc_hd__nand2_1 _26753_ (.A(_04633_),
    .B(_20637_),
    .Y(_04637_));
 sky130_fd_sc_hd__and2_1 _26754_ (.A(_04636_),
    .B(_04637_),
    .X(_02119_));
 sky130_fd_sc_hd__and3_1 _26755_ (.A(_18397_),
    .B(_04619_),
    .C(\irq_pending[25] ),
    .X(_04638_));
 sky130_fd_sc_hd__a221o_1 _26756_ (.A1(_04630_),
    .A2(\reg_next_pc[25] ),
    .B1(_04634_),
    .B2(_01536_),
    .C1(_04638_),
    .X(_02120_));
 sky130_fd_sc_hd__nor2_2 _26757_ (.A(_20643_),
    .B(_04636_),
    .Y(_04639_));
 sky130_fd_sc_hd__and2_1 _26758_ (.A(_04636_),
    .B(_20643_),
    .X(_04640_));
 sky130_fd_sc_hd__nor2_1 _26759_ (.A(_04639_),
    .B(_04640_),
    .Y(_02121_));
 sky130_fd_sc_hd__and3_1 _26760_ (.A(_18400_),
    .B(_04619_),
    .C(\irq_pending[26] ),
    .X(_04641_));
 sky130_fd_sc_hd__a221o_1 _26761_ (.A1(_04630_),
    .A2(\reg_next_pc[26] ),
    .B1(_04634_),
    .B2(_01539_),
    .C1(_04641_),
    .X(_02122_));
 sky130_fd_sc_hd__nor2_1 _26762_ (.A(\reg_pc[27] ),
    .B(_04639_),
    .Y(_04642_));
 sky130_fd_sc_hd__nand2_1 _26763_ (.A(_04639_),
    .B(\reg_pc[27] ),
    .Y(_04643_));
 sky130_vsdinv _26764_ (.A(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__nor2_1 _26765_ (.A(_04642_),
    .B(_04644_),
    .Y(_02123_));
 sky130_fd_sc_hd__and3_1 _26766_ (.A(_18402_),
    .B(_18529_),
    .C(\irq_pending[27] ),
    .X(_04645_));
 sky130_fd_sc_hd__a221o_1 _26767_ (.A1(_04630_),
    .A2(\reg_next_pc[27] ),
    .B1(_04634_),
    .B2(_01542_),
    .C1(_04645_),
    .X(_02124_));
 sky130_fd_sc_hd__nor2_2 _26768_ (.A(_20659_),
    .B(_04643_),
    .Y(_04646_));
 sky130_fd_sc_hd__nor2_1 _26769_ (.A(\reg_pc[28] ),
    .B(_04644_),
    .Y(_04647_));
 sky130_fd_sc_hd__nor2_1 _26770_ (.A(_04646_),
    .B(_04647_),
    .Y(_02125_));
 sky130_fd_sc_hd__and3_1 _26771_ (.A(_18435_),
    .B(_18529_),
    .C(\irq_pending[28] ),
    .X(_04648_));
 sky130_fd_sc_hd__a221o_1 _26772_ (.A1(_04630_),
    .A2(\reg_next_pc[28] ),
    .B1(_04634_),
    .B2(_01545_),
    .C1(_04648_),
    .X(_02126_));
 sky130_fd_sc_hd__nor2_1 _26773_ (.A(\reg_pc[29] ),
    .B(_04646_),
    .Y(_04649_));
 sky130_fd_sc_hd__and2_1 _26774_ (.A(_04646_),
    .B(\reg_pc[29] ),
    .X(_04650_));
 sky130_fd_sc_hd__nor2_1 _26775_ (.A(_04649_),
    .B(_04650_),
    .Y(_02127_));
 sky130_fd_sc_hd__and3_1 _26776_ (.A(_18343_),
    .B(_18485_),
    .C(_01548_),
    .X(_04651_));
 sky130_fd_sc_hd__a221o_1 _26777_ (.A1(_04581_),
    .A2(\reg_next_pc[29] ),
    .B1(_18437_),
    .B2(_18530_),
    .C1(_04651_),
    .X(_02128_));
 sky130_fd_sc_hd__or2_1 _26778_ (.A(\reg_pc[30] ),
    .B(_04650_),
    .X(_04652_));
 sky130_fd_sc_hd__nand2_1 _26779_ (.A(_04650_),
    .B(\reg_pc[30] ),
    .Y(_04653_));
 sky130_fd_sc_hd__and2_1 _26780_ (.A(_04652_),
    .B(_04653_),
    .X(_02129_));
 sky130_fd_sc_hd__and3_1 _26781_ (.A(_18434_),
    .B(_18529_),
    .C(\irq_pending[30] ),
    .X(_04654_));
 sky130_fd_sc_hd__a221o_1 _26782_ (.A1(_04581_),
    .A2(\reg_next_pc[30] ),
    .B1(_04634_),
    .B2(_01551_),
    .C1(_04654_),
    .X(_02130_));
 sky130_fd_sc_hd__xor2_1 _26783_ (.A(_20683_),
    .B(_04653_),
    .X(_02131_));
 sky130_fd_sc_hd__and3_1 _26784_ (.A(_18438_),
    .B(_18529_),
    .C(\irq_pending[31] ),
    .X(_04655_));
 sky130_fd_sc_hd__a221o_1 _26785_ (.A1(_04581_),
    .A2(\reg_next_pc[31] ),
    .B1(_04551_),
    .B2(_01554_),
    .C1(_04655_),
    .X(_02132_));
 sky130_fd_sc_hd__nor2_8 _26786_ (.A(instr_xor),
    .B(instr_xori),
    .Y(_04656_));
 sky130_vsdinv _26787_ (.A(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__nor2_4 _26788_ (.A(instr_sll),
    .B(instr_slli),
    .Y(_04658_));
 sky130_vsdinv _26789_ (.A(_04658_),
    .Y(_04659_));
 sky130_fd_sc_hd__clkbuf_2 _26790_ (.A(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__or3_2 _26791_ (.A(is_compare),
    .B(_04657_),
    .C(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_2 _26792_ (.A(_18506_),
    .X(_04662_));
 sky130_fd_sc_hd__buf_2 _26793_ (.A(_04662_),
    .X(_04663_));
 sky130_vsdinv _26794_ (.A(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__nor2_8 _26795_ (.A(instr_or),
    .B(instr_ori),
    .Y(_04665_));
 sky130_fd_sc_hd__clkbuf_2 _26796_ (.A(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__clkbuf_2 _26797_ (.A(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__nor2_8 _26798_ (.A(instr_and),
    .B(instr_andi),
    .Y(_04668_));
 sky130_fd_sc_hd__clkbuf_2 _26799_ (.A(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__and4b_4 _26800_ (.A_N(_04661_),
    .B(_04664_),
    .C(_04667_),
    .D(_04669_),
    .X(_02133_));
 sky130_fd_sc_hd__buf_2 _26801_ (.A(_04662_),
    .X(_04670_));
 sky130_fd_sc_hd__clkbuf_2 _26802_ (.A(_04657_),
    .X(_04671_));
 sky130_fd_sc_hd__clkbuf_2 _26803_ (.A(_04660_),
    .X(_04672_));
 sky130_vsdinv _26804_ (.A(_04668_),
    .Y(_04673_));
 sky130_fd_sc_hd__and3_1 _26805_ (.A(_04673_),
    .B(_19454_),
    .C(_19820_),
    .X(_04674_));
 sky130_vsdinv _26806_ (.A(_00343_),
    .Y(_04675_));
 sky130_vsdinv _26807_ (.A(_04665_),
    .Y(_04676_));
 sky130_fd_sc_hd__nand2_1 _26808_ (.A(_20202_),
    .B(_20119_),
    .Y(_04677_));
 sky130_fd_sc_hd__a22o_1 _26809_ (.A1(_04675_),
    .A2(is_compare),
    .B1(_04676_),
    .B2(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__a211o_1 _26810_ (.A1(\alu_shl[0] ),
    .A2(_04672_),
    .B1(_04674_),
    .C1(_04678_),
    .X(_04679_));
 sky130_fd_sc_hd__a221o_1 _26811_ (.A1(\alu_shr[0] ),
    .A2(_04670_),
    .B1(_02591_),
    .B2(_04671_),
    .C1(_04679_),
    .X(_02134_));
 sky130_fd_sc_hd__buf_2 _26812_ (.A(_04676_),
    .X(_04680_));
 sky130_fd_sc_hd__a2bb2o_1 _26813_ (.A1_N(_20340_),
    .A2_N(_04669_),
    .B1(\alu_shl[1] ),
    .B2(_04672_),
    .X(_04681_));
 sky130_fd_sc_hd__clkbuf_2 _26814_ (.A(_04656_),
    .X(_04682_));
 sky130_fd_sc_hd__clkbuf_2 _26815_ (.A(_04662_),
    .X(_04683_));
 sky130_fd_sc_hd__a2bb2o_1 _26816_ (.A1_N(_20341_),
    .A2_N(_04682_),
    .B1(\alu_shr[1] ),
    .B2(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__a211o_1 _26817_ (.A1(_20339_),
    .A2(_04680_),
    .B1(_04681_),
    .C1(_04684_),
    .X(_02135_));
 sky130_fd_sc_hd__buf_2 _26818_ (.A(_04673_),
    .X(_04685_));
 sky130_fd_sc_hd__and3_1 _26819_ (.A(_04685_),
    .B(net222),
    .C(_19817_),
    .X(_04686_));
 sky130_fd_sc_hd__clkbuf_2 _26820_ (.A(_04659_),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_2 _26821_ (.A(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__a2bb2o_1 _26822_ (.A1_N(_20287_),
    .A2_N(_04667_),
    .B1(\alu_shl[2] ),
    .B2(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__buf_2 _26823_ (.A(_04656_),
    .X(_04690_));
 sky130_fd_sc_hd__nor2_1 _26824_ (.A(_04690_),
    .B(_20290_),
    .Y(_04691_));
 sky130_fd_sc_hd__a2111o_1 _26825_ (.A1(\alu_shr[2] ),
    .A2(_04670_),
    .B1(_04686_),
    .C1(_04689_),
    .D1(_04691_),
    .X(_02136_));
 sky130_fd_sc_hd__buf_2 _26826_ (.A(_04662_),
    .X(_04692_));
 sky130_fd_sc_hd__nor2_1 _26827_ (.A(_20284_),
    .B(_20286_),
    .Y(_04693_));
 sky130_fd_sc_hd__buf_2 _26828_ (.A(_04673_),
    .X(_04694_));
 sky130_fd_sc_hd__buf_2 _26829_ (.A(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__buf_2 _26830_ (.A(_04665_),
    .X(_04696_));
 sky130_fd_sc_hd__a2bb2o_1 _26831_ (.A1_N(_20284_),
    .A2_N(_04696_),
    .B1(\alu_shl[3] ),
    .B2(_04660_),
    .X(_04697_));
 sky130_fd_sc_hd__a31o_1 _26832_ (.A1(net225),
    .A2(_19816_),
    .A3(_04695_),
    .B1(_04697_),
    .X(_04698_));
 sky130_fd_sc_hd__a221o_1 _26833_ (.A1(\alu_shr[3] ),
    .A2(_04692_),
    .B1(_04693_),
    .B2(_04671_),
    .C1(_04698_),
    .X(_02137_));
 sky130_fd_sc_hd__and3_1 _26834_ (.A(_04685_),
    .B(_19450_),
    .C(_19815_),
    .X(_04699_));
 sky130_fd_sc_hd__a2bb2o_1 _26835_ (.A1_N(_20276_),
    .A2_N(_04667_),
    .B1(\alu_shl[4] ),
    .B2(_04660_),
    .X(_04700_));
 sky130_fd_sc_hd__nor2_1 _26836_ (.A(_04690_),
    .B(_20279_),
    .Y(_04701_));
 sky130_fd_sc_hd__a2111o_1 _26837_ (.A1(\alu_shr[4] ),
    .A2(_04670_),
    .B1(_04699_),
    .C1(_04700_),
    .D1(_04701_),
    .X(_02138_));
 sky130_vsdinv _26838_ (.A(\alu_shr[5] ),
    .Y(_04702_));
 sky130_fd_sc_hd__clkbuf_2 _26839_ (.A(_04687_),
    .X(_04703_));
 sky130_fd_sc_hd__nand2_1 _26840_ (.A(_04703_),
    .B(\alu_shl[5] ),
    .Y(_04704_));
 sky130_fd_sc_hd__o221a_1 _26841_ (.A1(_20281_),
    .A2(_04668_),
    .B1(_20280_),
    .B2(_04667_),
    .C1(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__o221ai_1 _26842_ (.A1(_20282_),
    .A2(_04690_),
    .B1(_04702_),
    .B2(_04664_),
    .C1(_04705_),
    .Y(_02139_));
 sky130_fd_sc_hd__a2bb2o_1 _26843_ (.A1_N(_20330_),
    .A2_N(_04696_),
    .B1(\alu_shl[6] ),
    .B2(_04660_),
    .X(_04706_));
 sky130_fd_sc_hd__a31o_1 _26844_ (.A1(_19448_),
    .A2(_19813_),
    .A3(_04695_),
    .B1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__a221o_1 _26845_ (.A1(\alu_shr[6] ),
    .A2(_04692_),
    .B1(_20333_),
    .B2(_04671_),
    .C1(_04707_),
    .X(_02140_));
 sky130_fd_sc_hd__clkbuf_2 _26846_ (.A(_04666_),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_2 _26847_ (.A(_04659_),
    .X(_04709_));
 sky130_fd_sc_hd__a2bb2o_1 _26848_ (.A1_N(_20334_),
    .A2_N(_04708_),
    .B1(\alu_shl[7] ),
    .B2(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__a31o_1 _26849_ (.A1(net499),
    .A2(_19811_),
    .A3(_04695_),
    .B1(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__a221o_1 _26850_ (.A1(\alu_shr[7] ),
    .A2(_04692_),
    .B1(_20337_),
    .B2(_04671_),
    .C1(_04711_),
    .X(_02141_));
 sky130_fd_sc_hd__clkbuf_2 _26851_ (.A(_04694_),
    .X(_04712_));
 sky130_fd_sc_hd__a2bb2o_1 _26852_ (.A1_N(_20297_),
    .A2_N(_04708_),
    .B1(\alu_shl[8] ),
    .B2(_04709_),
    .X(_04713_));
 sky130_fd_sc_hd__a31o_1 _26853_ (.A1(_19445_),
    .A2(_19810_),
    .A3(_04712_),
    .B1(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__a221o_1 _26854_ (.A1(\alu_shr[8] ),
    .A2(_04692_),
    .B1(_20300_),
    .B2(_04671_),
    .C1(_04714_),
    .X(_02142_));
 sky130_fd_sc_hd__a2bb2o_1 _26855_ (.A1_N(_20307_),
    .A2_N(_04669_),
    .B1(\alu_shl[9] ),
    .B2(_04672_),
    .X(_04715_));
 sky130_fd_sc_hd__buf_2 _26856_ (.A(_04657_),
    .X(_04716_));
 sky130_fd_sc_hd__a22o_1 _26857_ (.A1(_20309_),
    .A2(_04716_),
    .B1(_04663_),
    .B2(\alu_shr[9] ),
    .X(_04717_));
 sky130_fd_sc_hd__a211o_1 _26858_ (.A1(_20306_),
    .A2(_04680_),
    .B1(_04715_),
    .C1(_04717_),
    .X(_02143_));
 sky130_fd_sc_hd__a2bb2o_1 _26859_ (.A1_N(_20293_),
    .A2_N(_04708_),
    .B1(\alu_shl[10] ),
    .B2(_04709_),
    .X(_04718_));
 sky130_fd_sc_hd__a31o_1 _26860_ (.A1(_19443_),
    .A2(_19808_),
    .A3(_04712_),
    .B1(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__a221o_1 _26861_ (.A1(\alu_shr[10] ),
    .A2(_04692_),
    .B1(_20296_),
    .B2(_04671_),
    .C1(_04719_),
    .X(_02144_));
 sky130_fd_sc_hd__clkbuf_2 _26862_ (.A(_04657_),
    .X(_04720_));
 sky130_fd_sc_hd__a2bb2o_1 _26863_ (.A1_N(_20301_),
    .A2_N(_04708_),
    .B1(\alu_shl[11] ),
    .B2(_04709_),
    .X(_04721_));
 sky130_fd_sc_hd__a31o_1 _26864_ (.A1(_19442_),
    .A2(_19807_),
    .A3(_04712_),
    .B1(_04721_),
    .X(_04722_));
 sky130_fd_sc_hd__a221o_1 _26865_ (.A1(\alu_shr[11] ),
    .A2(_04692_),
    .B1(_20304_),
    .B2(_04720_),
    .C1(_04722_),
    .X(_02145_));
 sky130_fd_sc_hd__and3_1 _26866_ (.A(_04694_),
    .B(_19441_),
    .C(_19806_),
    .X(_04723_));
 sky130_fd_sc_hd__a2bb2o_1 _26867_ (.A1_N(_20324_),
    .A2_N(_04667_),
    .B1(\alu_shl[12] ),
    .B2(_04660_),
    .X(_04724_));
 sky130_fd_sc_hd__nor2_1 _26868_ (.A(_04690_),
    .B(_20327_),
    .Y(_04725_));
 sky130_fd_sc_hd__a2111o_1 _26869_ (.A1(\alu_shr[12] ),
    .A2(_04670_),
    .B1(_04723_),
    .C1(_04724_),
    .D1(_04725_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_2 _26870_ (.A(_04662_),
    .X(_04726_));
 sky130_fd_sc_hd__a2bb2o_1 _26871_ (.A1_N(_20311_),
    .A2_N(_04708_),
    .B1(\alu_shl[13] ),
    .B2(_04709_),
    .X(_04727_));
 sky130_fd_sc_hd__a31o_1 _26872_ (.A1(_19440_),
    .A2(_19804_),
    .A3(_04712_),
    .B1(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__a221o_1 _26873_ (.A1(\alu_shr[13] ),
    .A2(_04726_),
    .B1(_20314_),
    .B2(_04720_),
    .C1(_04728_),
    .X(_02147_));
 sky130_fd_sc_hd__a2bb2o_1 _26874_ (.A1_N(_20317_),
    .A2_N(_04669_),
    .B1(\alu_shl[14] ),
    .B2(_04703_),
    .X(_04729_));
 sky130_fd_sc_hd__a22o_1 _26875_ (.A1(_20319_),
    .A2(_04657_),
    .B1(_04663_),
    .B2(\alu_shr[14] ),
    .X(_04730_));
 sky130_fd_sc_hd__a211o_1 _26876_ (.A1(_20316_),
    .A2(_04680_),
    .B1(_04729_),
    .C1(_04730_),
    .X(_02148_));
 sky130_vsdinv _26877_ (.A(_20320_),
    .Y(_04731_));
 sky130_fd_sc_hd__a22o_1 _26878_ (.A1(_04672_),
    .A2(\alu_shl[15] ),
    .B1(_20322_),
    .B2(_04695_),
    .X(_04732_));
 sky130_fd_sc_hd__a2bb2o_1 _26879_ (.A1_N(_04682_),
    .A2_N(_20323_),
    .B1(\alu_shr[15] ),
    .B2(_04683_),
    .X(_04733_));
 sky130_fd_sc_hd__a211o_1 _26880_ (.A1(_04731_),
    .A2(_04680_),
    .B1(_04732_),
    .C1(_04733_),
    .X(_02149_));
 sky130_fd_sc_hd__nor3_1 _26881_ (.A(_20261_),
    .B(_04690_),
    .C(_20263_),
    .Y(_04734_));
 sky130_fd_sc_hd__and3_1 _26882_ (.A(_04685_),
    .B(_19436_),
    .C(_19801_),
    .X(_04735_));
 sky130_fd_sc_hd__a2bb2o_1 _26883_ (.A1_N(_20261_),
    .A2_N(_04667_),
    .B1(\alu_shl[16] ),
    .B2(_04703_),
    .X(_04736_));
 sky130_fd_sc_hd__a2111o_2 _26884_ (.A1(_04670_),
    .A2(\alu_shr[16] ),
    .B1(_04734_),
    .C1(_04735_),
    .D1(_04736_),
    .X(_02150_));
 sky130_fd_sc_hd__a2bb2o_1 _26885_ (.A1_N(_20265_),
    .A2_N(_04708_),
    .B1(\alu_shl[17] ),
    .B2(_04709_),
    .X(_04737_));
 sky130_fd_sc_hd__a31o_1 _26886_ (.A1(net346),
    .A2(_19800_),
    .A3(_04712_),
    .B1(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__a221o_1 _26887_ (.A1(\alu_shr[17] ),
    .A2(_04726_),
    .B1(_20268_),
    .B2(_04720_),
    .C1(_04738_),
    .X(_02151_));
 sky130_fd_sc_hd__nor2_2 _26888_ (.A(_20258_),
    .B(_20260_),
    .Y(_04739_));
 sky130_fd_sc_hd__a2bb2o_1 _26889_ (.A1_N(_20258_),
    .A2_N(_04666_),
    .B1(\alu_shl[18] ),
    .B2(_04687_),
    .X(_04740_));
 sky130_fd_sc_hd__a31o_1 _26890_ (.A1(_19435_),
    .A2(_19799_),
    .A3(_04712_),
    .B1(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__a221o_1 _26891_ (.A1(\alu_shr[18] ),
    .A2(_04726_),
    .B1(_04739_),
    .B2(_04720_),
    .C1(_04741_),
    .X(_02152_));
 sky130_fd_sc_hd__a2bb2o_1 _26892_ (.A1_N(_20269_),
    .A2_N(_04666_),
    .B1(\alu_shl[19] ),
    .B2(_04687_),
    .X(_04742_));
 sky130_fd_sc_hd__a31o_1 _26893_ (.A1(net348),
    .A2(_19797_),
    .A3(_04685_),
    .B1(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__a221o_1 _26894_ (.A1(\alu_shr[19] ),
    .A2(_04726_),
    .B1(_20272_),
    .B2(_04720_),
    .C1(_04743_),
    .X(_02153_));
 sky130_fd_sc_hd__a2bb2o_1 _26895_ (.A1_N(_20246_),
    .A2_N(_04669_),
    .B1(\alu_shl[20] ),
    .B2(_04703_),
    .X(_04744_));
 sky130_fd_sc_hd__a2bb2o_1 _26896_ (.A1_N(_20247_),
    .A2_N(_04682_),
    .B1(\alu_shr[20] ),
    .B2(_04683_),
    .X(_04745_));
 sky130_fd_sc_hd__a211o_2 _26897_ (.A1(_20245_),
    .A2(_04680_),
    .B1(_04744_),
    .C1(_04745_),
    .X(_02154_));
 sky130_fd_sc_hd__a2bb2o_1 _26898_ (.A1_N(_20252_),
    .A2_N(_04666_),
    .B1(\alu_shl[21] ),
    .B2(_04687_),
    .X(_04746_));
 sky130_fd_sc_hd__a31o_1 _26899_ (.A1(_19433_),
    .A2(_19795_),
    .A3(_04685_),
    .B1(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__a221o_1 _26900_ (.A1(\alu_shr[21] ),
    .A2(_04726_),
    .B1(_20255_),
    .B2(_04720_),
    .C1(_04747_),
    .X(_02155_));
 sky130_fd_sc_hd__nor2_1 _26901_ (.A(_20241_),
    .B(_20243_),
    .Y(_04748_));
 sky130_fd_sc_hd__a2bb2o_1 _26902_ (.A1_N(_20241_),
    .A2_N(_04666_),
    .B1(\alu_shl[22] ),
    .B2(_04687_),
    .X(_04749_));
 sky130_fd_sc_hd__a31o_1 _26903_ (.A1(_19432_),
    .A2(_19794_),
    .A3(_04685_),
    .B1(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__a221o_2 _26904_ (.A1(\alu_shr[22] ),
    .A2(_04726_),
    .B1(_04748_),
    .B2(_04716_),
    .C1(_04750_),
    .X(_02156_));
 sky130_vsdinv _26905_ (.A(_20248_),
    .Y(_04751_));
 sky130_fd_sc_hd__a22o_1 _26906_ (.A1(_04672_),
    .A2(\alu_shl[23] ),
    .B1(_20250_),
    .B2(_04695_),
    .X(_04752_));
 sky130_fd_sc_hd__a2bb2o_1 _26907_ (.A1_N(_04682_),
    .A2_N(_20251_),
    .B1(\alu_shr[23] ),
    .B2(_04683_),
    .X(_04753_));
 sky130_fd_sc_hd__a211o_1 _26908_ (.A1(_04751_),
    .A2(_04680_),
    .B1(_04752_),
    .C1(_04753_),
    .X(_02157_));
 sky130_fd_sc_hd__a2bb2o_1 _26909_ (.A1_N(_20219_),
    .A2_N(_04669_),
    .B1(\alu_shl[24] ),
    .B2(_04703_),
    .X(_04754_));
 sky130_fd_sc_hd__a2bb2o_1 _26910_ (.A1_N(_20220_),
    .A2_N(_04682_),
    .B1(\alu_shr[24] ),
    .B2(_04683_),
    .X(_04755_));
 sky130_fd_sc_hd__a211o_1 _26911_ (.A1(_20218_),
    .A2(_04676_),
    .B1(_04754_),
    .C1(_04755_),
    .X(_02158_));
 sky130_fd_sc_hd__nor2_1 _26912_ (.A(_20204_),
    .B(_04696_),
    .Y(_04756_));
 sky130_fd_sc_hd__a221o_1 _26913_ (.A1(_04688_),
    .A2(\alu_shl[25] ),
    .B1(_20206_),
    .B2(_04694_),
    .C1(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__a221o_1 _26914_ (.A1(\alu_shr[25] ),
    .A2(_04663_),
    .B1(_20207_),
    .B2(_04716_),
    .C1(_04757_),
    .X(_02159_));
 sky130_vsdinv _26915_ (.A(_20209_),
    .Y(_04758_));
 sky130_fd_sc_hd__a22o_1 _26916_ (.A1(_04672_),
    .A2(\alu_shl[26] ),
    .B1(_20211_),
    .B2(_04695_),
    .X(_04759_));
 sky130_fd_sc_hd__a2bb2o_1 _26917_ (.A1_N(_04656_),
    .A2_N(_20212_),
    .B1(\alu_shr[26] ),
    .B2(_04683_),
    .X(_04760_));
 sky130_fd_sc_hd__a211o_1 _26918_ (.A1(_04758_),
    .A2(_04676_),
    .B1(_04759_),
    .C1(_04760_),
    .X(_02160_));
 sky130_vsdinv _26919_ (.A(_20216_),
    .Y(_04761_));
 sky130_fd_sc_hd__nor2_1 _26920_ (.A(_20215_),
    .B(_04668_),
    .Y(_04762_));
 sky130_fd_sc_hd__a221o_1 _26921_ (.A1(_04688_),
    .A2(\alu_shl[27] ),
    .B1(_20214_),
    .B2(_04676_),
    .C1(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__a221o_1 _26922_ (.A1(_04670_),
    .A2(\alu_shr[27] ),
    .B1(_04761_),
    .B2(_04716_),
    .C1(_04763_),
    .X(_02161_));
 sky130_fd_sc_hd__nor2_1 _26923_ (.A(_20235_),
    .B(_04696_),
    .Y(_04764_));
 sky130_fd_sc_hd__a221o_1 _26924_ (.A1(_04688_),
    .A2(\alu_shl[28] ),
    .B1(_20237_),
    .B2(_04694_),
    .C1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__a221o_1 _26925_ (.A1(\alu_shr[28] ),
    .A2(_04663_),
    .B1(_20238_),
    .B2(_04716_),
    .C1(_04765_),
    .X(_02162_));
 sky130_fd_sc_hd__nor2_1 _26926_ (.A(_20230_),
    .B(_04696_),
    .Y(_04766_));
 sky130_fd_sc_hd__a221o_1 _26927_ (.A1(_04688_),
    .A2(\alu_shl[29] ),
    .B1(_20232_),
    .B2(_04694_),
    .C1(_04766_),
    .X(_04767_));
 sky130_fd_sc_hd__a221o_1 _26928_ (.A1(\alu_shr[29] ),
    .A2(_04663_),
    .B1(_20233_),
    .B2(_04716_),
    .C1(_04767_),
    .X(_02163_));
 sky130_fd_sc_hd__a2bb2o_1 _26929_ (.A1_N(_20227_),
    .A2_N(_04668_),
    .B1(\alu_shl[30] ),
    .B2(_04703_),
    .X(_04768_));
 sky130_fd_sc_hd__a2bb2o_1 _26930_ (.A1_N(_20228_),
    .A2_N(_04682_),
    .B1(\alu_shr[30] ),
    .B2(_04662_),
    .X(_04769_));
 sky130_fd_sc_hd__a211o_1 _26931_ (.A1(_20226_),
    .A2(_04676_),
    .B1(_04768_),
    .C1(_04769_),
    .X(_02164_));
 sky130_vsdinv _26932_ (.A(\alu_shr[31] ),
    .Y(_04770_));
 sky130_fd_sc_hd__nand2_1 _26933_ (.A(_04688_),
    .B(\alu_shl[31] ),
    .Y(_04771_));
 sky130_fd_sc_hd__o221a_1 _26934_ (.A1(_20222_),
    .A2(_04696_),
    .B1(_20223_),
    .B2(_04668_),
    .C1(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__o221ai_2 _26935_ (.A1(_20224_),
    .A2(_04690_),
    .B1(_04770_),
    .B2(_04664_),
    .C1(_04772_),
    .Y(_02165_));
 sky130_fd_sc_hd__and3_1 _26936_ (.A(_00289_),
    .B(_18320_),
    .C(_20360_),
    .X(_02166_));
 sky130_vsdinv _26937_ (.A(_04116_),
    .Y(net233));
 sky130_fd_sc_hd__clkbuf_2 _26938_ (.A(\mem_wordsize[1] ),
    .X(_04773_));
 sky130_fd_sc_hd__a22o_1 _26939_ (.A1(_19445_),
    .A2(_04188_),
    .B1(_19454_),
    .B2(_04773_),
    .X(_02167_));
 sky130_fd_sc_hd__a22o_1 _26940_ (.A1(_19444_),
    .A2(_04188_),
    .B1(_19453_),
    .B2(_04773_),
    .X(_02168_));
 sky130_fd_sc_hd__clkbuf_2 _26941_ (.A(_04112_),
    .X(_04774_));
 sky130_fd_sc_hd__a22o_1 _26942_ (.A1(_19443_),
    .A2(_04774_),
    .B1(_19452_),
    .B2(_04773_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _26943_ (.A1(_19442_),
    .A2(_04774_),
    .B1(_19451_),
    .B2(_04773_),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_1 _26944_ (.A1(_19441_),
    .A2(_04774_),
    .B1(_19450_),
    .B2(_04773_),
    .X(_02171_));
 sky130_fd_sc_hd__a22o_1 _26945_ (.A1(_19440_),
    .A2(_04774_),
    .B1(_19449_),
    .B2(_04773_),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_1 _26946_ (.A1(_19438_),
    .A2(_04774_),
    .B1(_19448_),
    .B2(\mem_wordsize[1] ),
    .X(_02173_));
 sky130_fd_sc_hd__a22o_1 _26947_ (.A1(_19437_),
    .A2(_04774_),
    .B1(net499),
    .B2(\mem_wordsize[1] ),
    .X(_02174_));
 sky130_fd_sc_hd__nor2_1 _26948_ (.A(_20202_),
    .B(_04496_),
    .Y(_02175_));
 sky130_fd_sc_hd__clkbuf_2 _26949_ (.A(_04114_),
    .X(_04775_));
 sky130_fd_sc_hd__nor2_1 _26950_ (.A(_02318_),
    .B(_04775_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_2 _26951_ (.A(_02321_),
    .B(_04775_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _26952_ (.A(_02324_),
    .B(_04775_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _26953_ (.A(_02327_),
    .B(_04775_),
    .Y(_02179_));
 sky130_fd_sc_hd__inv_2 _26954_ (.A(_19449_),
    .Y(_02330_));
 sky130_fd_sc_hd__nor2_1 _26955_ (.A(_02330_),
    .B(_04775_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _26956_ (.A(_02333_),
    .B(_04775_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_1 _26957_ (.A(_02336_),
    .B(_04114_),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_8 _26958_ (.A(_20364_),
    .B(_18486_),
    .Y(_02183_));
 sky130_fd_sc_hd__or2_1 _26959_ (.A(\irq_pending[3] ),
    .B(net26),
    .X(_02214_));
 sky130_fd_sc_hd__and2_1 _26960_ (.A(_02214_),
    .B(\irq_mask[3] ),
    .X(_02215_));
 sky130_vsdinv _26961_ (.A(_01700_),
    .Y(_02217_));
 sky130_fd_sc_hd__or2_1 _26962_ (.A(\irq_pending[4] ),
    .B(net27),
    .X(_02218_));
 sky130_fd_sc_hd__and2_1 _26963_ (.A(_02218_),
    .B(\irq_mask[4] ),
    .X(_02219_));
 sky130_fd_sc_hd__or2_1 _26964_ (.A(\irq_pending[5] ),
    .B(net28),
    .X(_02221_));
 sky130_fd_sc_hd__and2_1 _26965_ (.A(_02221_),
    .B(\irq_mask[5] ),
    .X(_02222_));
 sky130_fd_sc_hd__or2_1 _26966_ (.A(\irq_pending[6] ),
    .B(net29),
    .X(_02224_));
 sky130_fd_sc_hd__and2_1 _26967_ (.A(_02224_),
    .B(\irq_mask[6] ),
    .X(_02225_));
 sky130_fd_sc_hd__or2_1 _26968_ (.A(\irq_pending[7] ),
    .B(net518),
    .X(_02227_));
 sky130_fd_sc_hd__and2_1 _26969_ (.A(_02227_),
    .B(\irq_mask[7] ),
    .X(_02228_));
 sky130_fd_sc_hd__or2_1 _26970_ (.A(\irq_pending[8] ),
    .B(net31),
    .X(_02230_));
 sky130_fd_sc_hd__and2_1 _26971_ (.A(_02230_),
    .B(\irq_mask[8] ),
    .X(_02231_));
 sky130_fd_sc_hd__or2_1 _26972_ (.A(\irq_pending[9] ),
    .B(net32),
    .X(_02233_));
 sky130_fd_sc_hd__and2_1 _26973_ (.A(_02233_),
    .B(\irq_mask[9] ),
    .X(_02234_));
 sky130_fd_sc_hd__or2_1 _26974_ (.A(\irq_pending[10] ),
    .B(net522),
    .X(_02236_));
 sky130_fd_sc_hd__and2_1 _26975_ (.A(_02236_),
    .B(\irq_mask[10] ),
    .X(_02237_));
 sky130_fd_sc_hd__or2_1 _26976_ (.A(\irq_pending[11] ),
    .B(net3),
    .X(_02239_));
 sky130_fd_sc_hd__and2_1 _26977_ (.A(_02239_),
    .B(\irq_mask[11] ),
    .X(_02240_));
 sky130_fd_sc_hd__or2_1 _26978_ (.A(\irq_pending[12] ),
    .B(net4),
    .X(_02242_));
 sky130_fd_sc_hd__and2_1 _26979_ (.A(_02242_),
    .B(\irq_mask[12] ),
    .X(_02243_));
 sky130_fd_sc_hd__or2_1 _26980_ (.A(\irq_pending[13] ),
    .B(net5),
    .X(_02245_));
 sky130_fd_sc_hd__and2_1 _26981_ (.A(_02245_),
    .B(\irq_mask[13] ),
    .X(_02246_));
 sky130_fd_sc_hd__or2_1 _26982_ (.A(\irq_pending[14] ),
    .B(net6),
    .X(_02248_));
 sky130_fd_sc_hd__and2_1 _26983_ (.A(_02248_),
    .B(\irq_mask[14] ),
    .X(_02249_));
 sky130_fd_sc_hd__or2_1 _26984_ (.A(\irq_pending[15] ),
    .B(net510),
    .X(_02251_));
 sky130_fd_sc_hd__and2_1 _26985_ (.A(_02251_),
    .B(\irq_mask[15] ),
    .X(_02252_));
 sky130_fd_sc_hd__or2_1 _26986_ (.A(\irq_pending[16] ),
    .B(net8),
    .X(_02254_));
 sky130_fd_sc_hd__and2_1 _26987_ (.A(_02254_),
    .B(\irq_mask[16] ),
    .X(_02255_));
 sky130_fd_sc_hd__or2_1 _26988_ (.A(\irq_pending[17] ),
    .B(net9),
    .X(_02257_));
 sky130_fd_sc_hd__and2_1 _26989_ (.A(_02257_),
    .B(\irq_mask[17] ),
    .X(_02258_));
 sky130_fd_sc_hd__or2_1 _26990_ (.A(\irq_pending[18] ),
    .B(net10),
    .X(_02260_));
 sky130_fd_sc_hd__and2_1 _26991_ (.A(_02260_),
    .B(\irq_mask[18] ),
    .X(_02261_));
 sky130_fd_sc_hd__or2_1 _26992_ (.A(\irq_pending[19] ),
    .B(net11),
    .X(_02263_));
 sky130_fd_sc_hd__and2_1 _26993_ (.A(_02263_),
    .B(\irq_mask[19] ),
    .X(_02264_));
 sky130_fd_sc_hd__or2_1 _26994_ (.A(\irq_pending[20] ),
    .B(net524),
    .X(_02266_));
 sky130_fd_sc_hd__and2_1 _26995_ (.A(_02266_),
    .B(\irq_mask[20] ),
    .X(_02267_));
 sky130_fd_sc_hd__or2_1 _26996_ (.A(\irq_pending[21] ),
    .B(net523),
    .X(_02269_));
 sky130_fd_sc_hd__and2_1 _26997_ (.A(_02269_),
    .B(\irq_mask[21] ),
    .X(_02270_));
 sky130_fd_sc_hd__or2_1 _26998_ (.A(\irq_pending[22] ),
    .B(net15),
    .X(_02272_));
 sky130_fd_sc_hd__and2_1 _26999_ (.A(_02272_),
    .B(\irq_mask[22] ),
    .X(_02273_));
 sky130_fd_sc_hd__or2_1 _27000_ (.A(\irq_pending[23] ),
    .B(net16),
    .X(_02275_));
 sky130_fd_sc_hd__and2_1 _27001_ (.A(_02275_),
    .B(\irq_mask[23] ),
    .X(_02276_));
 sky130_fd_sc_hd__or2_1 _27002_ (.A(\irq_pending[24] ),
    .B(net17),
    .X(_02278_));
 sky130_fd_sc_hd__and2_1 _27003_ (.A(_02278_),
    .B(\irq_mask[24] ),
    .X(_02279_));
 sky130_fd_sc_hd__or2_1 _27004_ (.A(\irq_pending[25] ),
    .B(net18),
    .X(_02281_));
 sky130_fd_sc_hd__and2_1 _27005_ (.A(_02281_),
    .B(\irq_mask[25] ),
    .X(_02282_));
 sky130_fd_sc_hd__or2_1 _27006_ (.A(\irq_pending[26] ),
    .B(net19),
    .X(_02284_));
 sky130_fd_sc_hd__and2_1 _27007_ (.A(_02284_),
    .B(\irq_mask[26] ),
    .X(_02285_));
 sky130_fd_sc_hd__or2_1 _27008_ (.A(\irq_pending[27] ),
    .B(net521),
    .X(_02287_));
 sky130_fd_sc_hd__and2_1 _27009_ (.A(_02287_),
    .B(\irq_mask[27] ),
    .X(_02288_));
 sky130_fd_sc_hd__or2_1 _27010_ (.A(\irq_pending[28] ),
    .B(net520),
    .X(_02290_));
 sky130_fd_sc_hd__and2_1 _27011_ (.A(_02290_),
    .B(\irq_mask[28] ),
    .X(_02291_));
 sky130_fd_sc_hd__or2_1 _27012_ (.A(\irq_pending[29] ),
    .B(net22),
    .X(_02293_));
 sky130_fd_sc_hd__and2_1 _27013_ (.A(_02293_),
    .B(\irq_mask[29] ),
    .X(_02294_));
 sky130_fd_sc_hd__or2_1 _27014_ (.A(\irq_pending[30] ),
    .B(net24),
    .X(_02296_));
 sky130_fd_sc_hd__and2_1 _27015_ (.A(_02296_),
    .B(\irq_mask[30] ),
    .X(_02297_));
 sky130_fd_sc_hd__or2_1 _27016_ (.A(\irq_pending[31] ),
    .B(net519),
    .X(_02299_));
 sky130_fd_sc_hd__and2_1 _27017_ (.A(_02299_),
    .B(\irq_mask[31] ),
    .X(_02300_));
 sky130_fd_sc_hd__or4_4 _27018_ (.A(\timer[7] ),
    .B(\timer[6] ),
    .C(\timer[17] ),
    .D(\timer[19] ),
    .X(_04776_));
 sky130_fd_sc_hd__or4_4 _27019_ (.A(\timer[1] ),
    .B(\timer[3] ),
    .C(\timer[2] ),
    .D(_20368_),
    .X(_04777_));
 sky130_fd_sc_hd__nor2_1 _27020_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__and3_1 _27021_ (.A(_20395_),
    .B(_04498_),
    .C(_04484_),
    .X(_04779_));
 sky130_fd_sc_hd__and3_1 _27022_ (.A(_04779_),
    .B(_20402_),
    .C(_20385_),
    .X(_04780_));
 sky130_fd_sc_hd__and3_1 _27023_ (.A(_04380_),
    .B(_04422_),
    .C(_20390_),
    .X(_04781_));
 sky130_fd_sc_hd__and4_1 _27024_ (.A(_04781_),
    .B(_20379_),
    .C(_04273_),
    .D(_20380_),
    .X(_04782_));
 sky130_fd_sc_hd__nor2_1 _27025_ (.A(\timer[23] ),
    .B(\timer[22] ),
    .Y(_04783_));
 sky130_fd_sc_hd__and3_1 _27026_ (.A(_04783_),
    .B(_20365_),
    .C(_20376_),
    .X(_04784_));
 sky130_fd_sc_hd__a41o_1 _27027_ (.A1(_04778_),
    .A2(_04780_),
    .A3(_04782_),
    .A4(_04784_),
    .B1(\irq_pending[0] ),
    .X(_02302_));
 sky130_fd_sc_hd__or2_1 _27028_ (.A(_02303_),
    .B(net1),
    .X(_02304_));
 sky130_fd_sc_hd__and2_1 _27029_ (.A(_02304_),
    .B(\irq_mask[0] ),
    .X(_02305_));
 sky130_fd_sc_hd__nor2_2 _27030_ (.A(\irq_pending[2] ),
    .B(net23),
    .Y(_02307_));
 sky130_fd_sc_hd__or2_1 _27031_ (.A(_18623_),
    .B(_02307_),
    .X(_02308_));
 sky130_fd_sc_hd__nor2_1 _27032_ (.A(_02310_),
    .B(_18589_),
    .Y(_02311_));
 sky130_fd_sc_hd__or2_1 _27033_ (.A(_20134_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__or2_1 _27034_ (.A(_02313_),
    .B(_20134_),
    .X(_02314_));
 sky130_fd_sc_hd__or2_1 _27035_ (.A(_02316_),
    .B(_20134_),
    .X(_02317_));
 sky130_fd_sc_hd__nor2_1 _27036_ (.A(_19803_),
    .B(_02357_),
    .Y(_04785_));
 sky130_fd_sc_hd__or3_1 _27037_ (.A(_02351_),
    .B(_19806_),
    .C(_20314_),
    .X(_04786_));
 sky130_fd_sc_hd__nand2_1 _27038_ (.A(_20312_),
    .B(_19440_),
    .Y(_04787_));
 sky130_fd_sc_hd__a21oi_1 _27039_ (.A1(_04786_),
    .A2(_04787_),
    .B1(_20319_),
    .Y(_04788_));
 sky130_fd_sc_hd__o21ai_1 _27040_ (.A1(_04785_),
    .A2(_04788_),
    .B1(_20323_),
    .Y(_04789_));
 sky130_vsdinv _27041_ (.A(_20120_),
    .Y(_04790_));
 sky130_fd_sc_hd__nor2_2 _27042_ (.A(_20118_),
    .B(_04790_),
    .Y(_00049_));
 sky130_fd_sc_hd__o21a_1 _27043_ (.A1(_20117_),
    .A2(_00048_),
    .B1(_19818_),
    .X(_04791_));
 sky130_fd_sc_hd__nand2_1 _27044_ (.A(_20285_),
    .B(net225),
    .Y(_04792_));
 sky130_fd_sc_hd__or3_2 _27045_ (.A(_20116_),
    .B(_19817_),
    .C(_04693_),
    .X(_04793_));
 sky130_fd_sc_hd__o311a_1 _27046_ (.A1(_00049_),
    .A2(_04791_),
    .A3(_20291_),
    .B1(_04792_),
    .C1(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__or2_1 _27047_ (.A(_20283_),
    .B(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__or2_1 _27048_ (.A(_19814_),
    .B(_02330_),
    .X(_04796_));
 sky130_fd_sc_hd__or3b_2 _27049_ (.A(_20110_),
    .B(_19815_),
    .C_N(_20282_),
    .X(_04797_));
 sky130_fd_sc_hd__a31o_1 _27050_ (.A1(_04795_),
    .A2(_04796_),
    .A3(_04797_),
    .B1(_20333_),
    .X(_04798_));
 sky130_fd_sc_hd__nand2_1 _27051_ (.A(_20331_),
    .B(net228),
    .Y(_04799_));
 sky130_fd_sc_hd__a21o_1 _27052_ (.A1(_04798_),
    .A2(_04799_),
    .B1(_20337_),
    .X(_04800_));
 sky130_fd_sc_hd__nand2_1 _27053_ (.A(_20335_),
    .B(net229),
    .Y(_04801_));
 sky130_fd_sc_hd__a21o_1 _27054_ (.A1(_04800_),
    .A2(_04801_),
    .B1(_20310_),
    .X(_04802_));
 sky130_fd_sc_hd__nand2_1 _27055_ (.A(_20302_),
    .B(_19442_),
    .Y(_04803_));
 sky130_fd_sc_hd__and3_1 _27056_ (.A(_20308_),
    .B(_19445_),
    .C(_20298_),
    .X(_04804_));
 sky130_fd_sc_hd__a21oi_1 _27057_ (.A1(_19444_),
    .A2(_20305_),
    .B1(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__or2_1 _27058_ (.A(_20296_),
    .B(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__nand2_1 _27059_ (.A(_20294_),
    .B(_19443_),
    .Y(_04807_));
 sky130_fd_sc_hd__a21o_1 _27060_ (.A1(_04806_),
    .A2(_04807_),
    .B1(_20304_),
    .X(_04808_));
 sky130_fd_sc_hd__a31o_1 _27061_ (.A1(_04802_),
    .A2(_04803_),
    .A3(_04808_),
    .B1(_20329_),
    .X(_04809_));
 sky130_fd_sc_hd__o211a_1 _27062_ (.A1(_02360_),
    .A2(_19802_),
    .B1(_04789_),
    .C1(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__inv_2 _27063_ (.A(_19429_),
    .Y(_02396_));
 sky130_fd_sc_hd__nor2_1 _27064_ (.A(_19790_),
    .B(_02390_),
    .Y(_04811_));
 sky130_fd_sc_hd__and3_1 _27065_ (.A(_20208_),
    .B(net354),
    .C(_20217_),
    .X(_04812_));
 sky130_fd_sc_hd__o21ai_1 _27066_ (.A1(_04811_),
    .A2(_04812_),
    .B1(_20212_),
    .Y(_04813_));
 sky130_fd_sc_hd__nand2_1 _27067_ (.A(_20210_),
    .B(net356),
    .Y(_04814_));
 sky130_fd_sc_hd__a21o_1 _27068_ (.A1(_04813_),
    .A2(_04814_),
    .B1(_04761_),
    .X(_04815_));
 sky130_fd_sc_hd__o21ai_1 _27069_ (.A1(_02396_),
    .A2(_19789_),
    .B1(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__nor2_1 _27070_ (.A(_19788_),
    .B(_02402_),
    .Y(_04817_));
 sky130_fd_sc_hd__a31o_1 _27071_ (.A1(_04816_),
    .A2(_20234_),
    .A3(_20239_),
    .B1(_04817_),
    .X(_04818_));
 sky130_fd_sc_hd__a31o_1 _27072_ (.A1(net358),
    .A2(_20236_),
    .A3(_20234_),
    .B1(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__nand2_1 _27073_ (.A(_04819_),
    .B(_20229_),
    .Y(_04820_));
 sky130_fd_sc_hd__or3_1 _27074_ (.A(_02363_),
    .B(_19801_),
    .C(_20268_),
    .X(_04821_));
 sky130_fd_sc_hd__nand2_1 _27075_ (.A(_20266_),
    .B(net346),
    .Y(_04822_));
 sky130_fd_sc_hd__a21o_1 _27076_ (.A1(_04821_),
    .A2(_04822_),
    .B1(_04739_),
    .X(_04823_));
 sky130_fd_sc_hd__nand2_1 _27077_ (.A(_20259_),
    .B(_19435_),
    .Y(_04824_));
 sky130_fd_sc_hd__a21o_1 _27078_ (.A1(_04823_),
    .A2(_04824_),
    .B1(_20272_),
    .X(_04825_));
 sky130_fd_sc_hd__o21ai_1 _27079_ (.A1(_02372_),
    .A2(_19797_),
    .B1(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__nor2_1 _27080_ (.A(_19794_),
    .B(_02381_),
    .Y(_04827_));
 sky130_fd_sc_hd__nand2_1 _27081_ (.A(_20253_),
    .B(_19433_),
    .Y(_04828_));
 sky130_fd_sc_hd__o31a_1 _27082_ (.A1(_02375_),
    .A2(_19796_),
    .A3(_20255_),
    .B1(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__nor2_1 _27083_ (.A(_04748_),
    .B(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__o21a_1 _27084_ (.A1(_04827_),
    .A2(_04830_),
    .B1(_20251_),
    .X(_04831_));
 sky130_fd_sc_hd__a221o_1 _27085_ (.A1(_19431_),
    .A2(_20249_),
    .B1(_04826_),
    .B2(_20257_),
    .C1(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__and3_1 _27086_ (.A(_20224_),
    .B(_19428_),
    .C(_20225_),
    .X(_04833_));
 sky130_fd_sc_hd__a21oi_1 _27087_ (.A1(_04832_),
    .A2(_20240_),
    .B1(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__o211a_1 _27088_ (.A1(_20275_),
    .A2(_04810_),
    .B1(_04820_),
    .C1(_04834_),
    .X(_04835_));
 sky130_fd_sc_hd__nand2_2 _27089_ (.A(_20684_),
    .B(_18471_),
    .Y(_04836_));
 sky130_fd_sc_hd__a21oi_4 _27090_ (.A1(_04835_),
    .A2(_04836_),
    .B1(_00000_),
    .Y(_00002_));
 sky130_fd_sc_hd__nand2_1 _27091_ (.A(_04835_),
    .B(_20224_),
    .Y(_04837_));
 sky130_fd_sc_hd__o211a_1 _27092_ (.A1(_20343_),
    .A2(_20275_),
    .B1(_04836_),
    .C1(_04837_),
    .X(_00001_));
 sky130_vsdinv _27093_ (.A(\pcpi_mul.rs2[0] ),
    .Y(_04838_));
 sky130_fd_sc_hd__clkbuf_4 _27094_ (.A(_04838_),
    .X(_04839_));
 sky130_vsdinv _27095_ (.A(_19932_),
    .Y(_04840_));
 sky130_fd_sc_hd__clkbuf_2 _27096_ (.A(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__clkbuf_8 _27097_ (.A(net453),
    .X(_04842_));
 sky130_fd_sc_hd__nor2_2 _27098_ (.A(_04839_),
    .B(_04842_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand2_1 _27099_ (.A(_19453_),
    .B(_19454_),
    .Y(_04843_));
 sky130_fd_sc_hd__nand2_1 _27100_ (.A(_04790_),
    .B(_04843_),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_1 _27101_ (.A(_19818_),
    .B(_02320_),
    .Y(_04844_));
 sky130_fd_sc_hd__nand2_1 _27102_ (.A(_19818_),
    .B(_02320_),
    .Y(_04845_));
 sky130_fd_sc_hd__or2b_1 _27103_ (.A(_04844_),
    .B_N(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__xor2_1 _27104_ (.A(_20203_),
    .B(_04846_),
    .X(_02602_));
 sky130_vsdinv _27105_ (.A(_20121_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _27106_ (.A(_04790_),
    .B(_19452_),
    .Y(_04848_));
 sky130_fd_sc_hd__nand2_1 _27107_ (.A(_04847_),
    .B(_04848_),
    .Y(_02322_));
 sky130_fd_sc_hd__or2_1 _27108_ (.A(net328),
    .B(_02323_),
    .X(_04849_));
 sky130_fd_sc_hd__nand2_1 _27109_ (.A(net328),
    .B(_02323_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand2_1 _27110_ (.A(_04849_),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__o21ai_2 _27111_ (.A1(_04844_),
    .A2(_20203_),
    .B1(_04845_),
    .Y(_04852_));
 sky130_fd_sc_hd__xnor2_1 _27112_ (.A(_04851_),
    .B(_04852_),
    .Y(_02613_));
 sky130_fd_sc_hd__nand2_1 _27113_ (.A(_04847_),
    .B(_19451_),
    .Y(_04853_));
 sky130_fd_sc_hd__nand2_1 _27114_ (.A(_04853_),
    .B(_20122_),
    .Y(_02325_));
 sky130_fd_sc_hd__nor2_1 _27115_ (.A(net331),
    .B(_02326_),
    .Y(_04854_));
 sky130_fd_sc_hd__nand2_1 _27116_ (.A(net331),
    .B(_02326_),
    .Y(_04855_));
 sky130_vsdinv _27117_ (.A(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__or2_1 _27118_ (.A(_04854_),
    .B(_04856_),
    .X(_04857_));
 sky130_fd_sc_hd__nand2_1 _27119_ (.A(_04852_),
    .B(_04849_),
    .Y(_04858_));
 sky130_fd_sc_hd__and2_1 _27120_ (.A(_04858_),
    .B(_04850_),
    .X(_04859_));
 sky130_fd_sc_hd__xor2_1 _27121_ (.A(_04857_),
    .B(_04859_),
    .X(_02616_));
 sky130_fd_sc_hd__or2_1 _27122_ (.A(net226),
    .B(_20122_),
    .X(_04860_));
 sky130_fd_sc_hd__nand2_1 _27123_ (.A(_20122_),
    .B(_19450_),
    .Y(_04861_));
 sky130_fd_sc_hd__nand2_1 _27124_ (.A(_04860_),
    .B(_04861_),
    .Y(_02328_));
 sky130_vsdinv _27125_ (.A(_02329_),
    .Y(_04862_));
 sky130_fd_sc_hd__nor2_1 _27126_ (.A(_20277_),
    .B(_04862_),
    .Y(_04863_));
 sky130_vsdinv _27127_ (.A(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__nor2_1 _27128_ (.A(net332),
    .B(_02329_),
    .Y(_04865_));
 sky130_vsdinv _27129_ (.A(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__nand2_1 _27130_ (.A(_04864_),
    .B(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__a21oi_2 _27131_ (.A1(_04858_),
    .A2(_04850_),
    .B1(_04854_),
    .Y(_04868_));
 sky130_fd_sc_hd__nor2_1 _27132_ (.A(_04856_),
    .B(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__xor2_1 _27133_ (.A(_04867_),
    .B(_04869_),
    .X(_02617_));
 sky130_fd_sc_hd__or2_1 _27134_ (.A(net227),
    .B(_04860_),
    .X(_04870_));
 sky130_fd_sc_hd__nand2_1 _27135_ (.A(_04860_),
    .B(_19449_),
    .Y(_04871_));
 sky130_fd_sc_hd__nand2_1 _27136_ (.A(_04870_),
    .B(_04871_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_1 _27137_ (.A(net333),
    .B(_02332_),
    .Y(_04872_));
 sky130_fd_sc_hd__nand2_1 _27138_ (.A(net333),
    .B(_02332_),
    .Y(_04873_));
 sky130_vsdinv _27139_ (.A(_04873_),
    .Y(_04874_));
 sky130_fd_sc_hd__or2_1 _27140_ (.A(_04872_),
    .B(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__o21ai_1 _27141_ (.A1(_04856_),
    .A2(_04868_),
    .B1(_04866_),
    .Y(_04876_));
 sky130_fd_sc_hd__and2_1 _27142_ (.A(_04876_),
    .B(_04864_),
    .X(_04877_));
 sky130_fd_sc_hd__xor2_1 _27143_ (.A(_04875_),
    .B(_04877_),
    .X(_02618_));
 sky130_fd_sc_hd__or2_1 _27144_ (.A(net228),
    .B(_04870_),
    .X(_04878_));
 sky130_fd_sc_hd__nand2_1 _27145_ (.A(_04870_),
    .B(_19448_),
    .Y(_04879_));
 sky130_fd_sc_hd__nand2_1 _27146_ (.A(_04878_),
    .B(_04879_),
    .Y(_02334_));
 sky130_fd_sc_hd__xor2_2 _27147_ (.A(net334),
    .B(_02335_),
    .X(_04880_));
 sky130_fd_sc_hd__a21oi_2 _27148_ (.A1(_04876_),
    .A2(_04864_),
    .B1(_04872_),
    .Y(_04881_));
 sky130_fd_sc_hd__or2_1 _27149_ (.A(_04874_),
    .B(_04881_),
    .X(_04882_));
 sky130_fd_sc_hd__or2_1 _27150_ (.A(_04880_),
    .B(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__nand2_1 _27151_ (.A(_04882_),
    .B(_04880_),
    .Y(_04884_));
 sky130_fd_sc_hd__and2_1 _27152_ (.A(_04883_),
    .B(_04884_),
    .X(_02619_));
 sky130_fd_sc_hd__nor2_1 _27153_ (.A(net229),
    .B(_04878_),
    .Y(_04885_));
 sky130_fd_sc_hd__and2_1 _27154_ (.A(_04878_),
    .B(net499),
    .X(_04886_));
 sky130_fd_sc_hd__or2_1 _27155_ (.A(_04885_),
    .B(_04886_),
    .X(_02337_));
 sky130_fd_sc_hd__nor2_1 _27156_ (.A(_19811_),
    .B(_02338_),
    .Y(_04887_));
 sky130_fd_sc_hd__and2_1 _27157_ (.A(net335),
    .B(_02338_),
    .X(_04888_));
 sky130_fd_sc_hd__nor2_1 _27158_ (.A(_04887_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__a21bo_1 _27159_ (.A1(_19813_),
    .A2(_02335_),
    .B1_N(_04884_),
    .X(_04890_));
 sky130_fd_sc_hd__xor2_1 _27160_ (.A(_04889_),
    .B(_04890_),
    .X(_02620_));
 sky130_fd_sc_hd__or2_1 _27161_ (.A(_02339_),
    .B(_04885_),
    .X(_04891_));
 sky130_fd_sc_hd__nand2_1 _27162_ (.A(_04885_),
    .B(_02339_),
    .Y(_04892_));
 sky130_fd_sc_hd__nand2_1 _27163_ (.A(_04891_),
    .B(_04892_),
    .Y(_02340_));
 sky130_fd_sc_hd__or2_1 _27164_ (.A(net336),
    .B(_02341_),
    .X(_04893_));
 sky130_fd_sc_hd__nand2_1 _27165_ (.A(_19810_),
    .B(_02341_),
    .Y(_04894_));
 sky130_fd_sc_hd__and2_1 _27166_ (.A(_04893_),
    .B(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__and2_1 _27167_ (.A(_04880_),
    .B(_04889_),
    .X(_04896_));
 sky130_fd_sc_hd__o21ai_2 _27168_ (.A1(_04874_),
    .A2(_04881_),
    .B1(_04896_),
    .Y(_04897_));
 sky130_vsdinv _27169_ (.A(_04887_),
    .Y(_04898_));
 sky130_fd_sc_hd__a31oi_4 _27170_ (.A1(_04898_),
    .A2(_19813_),
    .A3(_02335_),
    .B1(_04888_),
    .Y(_04899_));
 sky130_fd_sc_hd__nand2_1 _27171_ (.A(_04897_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__or2_1 _27172_ (.A(_04895_),
    .B(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__nand2_1 _27173_ (.A(_04900_),
    .B(_04895_),
    .Y(_04902_));
 sky130_fd_sc_hd__and2_1 _27174_ (.A(_04901_),
    .B(_04902_),
    .X(_02621_));
 sky130_fd_sc_hd__or2_1 _27175_ (.A(net369),
    .B(_04892_),
    .X(_04903_));
 sky130_fd_sc_hd__nand2_1 _27176_ (.A(_04892_),
    .B(_19444_),
    .Y(_04904_));
 sky130_fd_sc_hd__nand2_1 _27177_ (.A(_04903_),
    .B(_04904_),
    .Y(_02343_));
 sky130_fd_sc_hd__nor2_1 _27178_ (.A(_19809_),
    .B(_02344_),
    .Y(_04905_));
 sky130_fd_sc_hd__and2_1 _27179_ (.A(_19809_),
    .B(_02344_),
    .X(_04906_));
 sky130_fd_sc_hd__nor2_2 _27180_ (.A(_04905_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__nand2_1 _27181_ (.A(_04902_),
    .B(_04894_),
    .Y(_04908_));
 sky130_fd_sc_hd__xor2_1 _27182_ (.A(_04907_),
    .B(_04908_),
    .X(_02622_));
 sky130_fd_sc_hd__or2_1 _27183_ (.A(net339),
    .B(_04903_),
    .X(_04909_));
 sky130_fd_sc_hd__nand2_1 _27184_ (.A(_04903_),
    .B(_19443_),
    .Y(_04910_));
 sky130_fd_sc_hd__nand2_1 _27185_ (.A(_04909_),
    .B(_04910_),
    .Y(_02346_));
 sky130_fd_sc_hd__or2_1 _27186_ (.A(net307),
    .B(_02347_),
    .X(_04911_));
 sky130_fd_sc_hd__nand2_1 _27187_ (.A(_19808_),
    .B(_02347_),
    .Y(_04912_));
 sky130_fd_sc_hd__and2_1 _27188_ (.A(_04911_),
    .B(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__o21bai_1 _27189_ (.A1(_04894_),
    .A2(_04905_),
    .B1_N(_04906_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand2_1 _27190_ (.A(_04895_),
    .B(_04907_),
    .Y(_04915_));
 sky130_fd_sc_hd__a21oi_2 _27191_ (.A1(_04897_),
    .A2(_04899_),
    .B1(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__or3_2 _27192_ (.A(_04913_),
    .B(_04914_),
    .C(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__o21ai_2 _27193_ (.A1(_04914_),
    .A2(_04916_),
    .B1(_04913_),
    .Y(_04918_));
 sky130_fd_sc_hd__and2_1 _27194_ (.A(_04917_),
    .B(_04918_),
    .X(_02592_));
 sky130_fd_sc_hd__or2_1 _27195_ (.A(net340),
    .B(_04909_),
    .X(_04919_));
 sky130_fd_sc_hd__nand2_1 _27196_ (.A(_04909_),
    .B(_19442_),
    .Y(_04920_));
 sky130_fd_sc_hd__nand2_1 _27197_ (.A(_04919_),
    .B(_04920_),
    .Y(_02349_));
 sky130_fd_sc_hd__or2_1 _27198_ (.A(net308),
    .B(_02350_),
    .X(_04921_));
 sky130_fd_sc_hd__nand2_1 _27199_ (.A(_19807_),
    .B(_02350_),
    .Y(_04922_));
 sky130_fd_sc_hd__nand2_1 _27200_ (.A(_04921_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__a21oi_2 _27201_ (.A1(_04918_),
    .A2(_04912_),
    .B1(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__and3_1 _27202_ (.A(_04918_),
    .B(_04912_),
    .C(_04923_),
    .X(_04925_));
 sky130_fd_sc_hd__nor2_1 _27203_ (.A(_04924_),
    .B(_04925_),
    .Y(_02593_));
 sky130_fd_sc_hd__nor2_1 _27204_ (.A(net341),
    .B(_04919_),
    .Y(_04926_));
 sky130_fd_sc_hd__and2_1 _27205_ (.A(_04919_),
    .B(_19441_),
    .X(_04927_));
 sky130_fd_sc_hd__or2_1 _27206_ (.A(_04926_),
    .B(_04927_),
    .X(_02352_));
 sky130_vsdinv _27207_ (.A(_04922_),
    .Y(_04928_));
 sky130_fd_sc_hd__or2_1 _27208_ (.A(net309),
    .B(_02353_),
    .X(_04929_));
 sky130_fd_sc_hd__nand2_1 _27209_ (.A(_19806_),
    .B(_02353_),
    .Y(_04930_));
 sky130_fd_sc_hd__and2_1 _27210_ (.A(_04929_),
    .B(_04930_),
    .X(_04931_));
 sky130_fd_sc_hd__or3_2 _27211_ (.A(_04928_),
    .B(_04931_),
    .C(_04924_),
    .X(_04932_));
 sky130_fd_sc_hd__o21ai_2 _27212_ (.A1(_04928_),
    .A2(_04924_),
    .B1(_04931_),
    .Y(_04933_));
 sky130_fd_sc_hd__and2_1 _27213_ (.A(_04932_),
    .B(_04933_),
    .X(_02594_));
 sky130_fd_sc_hd__or2_1 _27214_ (.A(_02354_),
    .B(_04926_),
    .X(_04934_));
 sky130_fd_sc_hd__nand2_1 _27215_ (.A(_04926_),
    .B(_02354_),
    .Y(_04935_));
 sky130_fd_sc_hd__nand2_1 _27216_ (.A(_04934_),
    .B(_04935_),
    .Y(_02355_));
 sky130_fd_sc_hd__or2_1 _27217_ (.A(net310),
    .B(_02356_),
    .X(_04936_));
 sky130_fd_sc_hd__nand2_1 _27218_ (.A(_19804_),
    .B(_02356_),
    .Y(_04937_));
 sky130_fd_sc_hd__nand2_1 _27219_ (.A(_04936_),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21oi_2 _27220_ (.A1(_04933_),
    .A2(_04930_),
    .B1(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__and3_1 _27221_ (.A(_04933_),
    .B(_04930_),
    .C(_04938_),
    .X(_04940_));
 sky130_fd_sc_hd__nor2_1 _27222_ (.A(_04939_),
    .B(_04940_),
    .Y(_02595_));
 sky130_fd_sc_hd__or2_1 _27223_ (.A(net343),
    .B(_04935_),
    .X(_04941_));
 sky130_fd_sc_hd__nand2_1 _27224_ (.A(_04935_),
    .B(_19438_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2_1 _27225_ (.A(_04941_),
    .B(_04942_),
    .Y(_02358_));
 sky130_vsdinv _27226_ (.A(_04937_),
    .Y(_04943_));
 sky130_fd_sc_hd__or2_1 _27227_ (.A(net311),
    .B(_02359_),
    .X(_04944_));
 sky130_fd_sc_hd__nand2_1 _27228_ (.A(_19803_),
    .B(_02359_),
    .Y(_04945_));
 sky130_fd_sc_hd__and2_1 _27229_ (.A(_04944_),
    .B(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__or3_2 _27230_ (.A(_04943_),
    .B(_04946_),
    .C(_04939_),
    .X(_04947_));
 sky130_fd_sc_hd__o21ai_2 _27231_ (.A1(_04943_),
    .A2(_04939_),
    .B1(_04946_),
    .Y(_04948_));
 sky130_fd_sc_hd__and2_1 _27232_ (.A(_04947_),
    .B(_04948_),
    .X(_02596_));
 sky130_fd_sc_hd__or2_1 _27233_ (.A(net344),
    .B(_04941_),
    .X(_04949_));
 sky130_fd_sc_hd__nand2_1 _27234_ (.A(_04941_),
    .B(_19437_),
    .Y(_04950_));
 sky130_fd_sc_hd__nand2_1 _27235_ (.A(_04949_),
    .B(_04950_),
    .Y(_02361_));
 sky130_fd_sc_hd__or2_1 _27236_ (.A(net312),
    .B(_02362_),
    .X(_04951_));
 sky130_fd_sc_hd__nand2_1 _27237_ (.A(_19802_),
    .B(_02362_),
    .Y(_04952_));
 sky130_fd_sc_hd__nand2_1 _27238_ (.A(_04951_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__a21oi_2 _27239_ (.A1(_04948_),
    .A2(_04945_),
    .B1(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__and3_1 _27240_ (.A(_04948_),
    .B(_04945_),
    .C(_04953_),
    .X(_04955_));
 sky130_fd_sc_hd__nor2_1 _27241_ (.A(_04954_),
    .B(_04955_),
    .Y(_02597_));
 sky130_fd_sc_hd__nor2_1 _27242_ (.A(net345),
    .B(_04949_),
    .Y(_04956_));
 sky130_fd_sc_hd__and2_1 _27243_ (.A(_04949_),
    .B(_19436_),
    .X(_04957_));
 sky130_fd_sc_hd__or2_1 _27244_ (.A(_04956_),
    .B(_04957_),
    .X(_02364_));
 sky130_fd_sc_hd__xor2_1 _27245_ (.A(net313),
    .B(_02365_),
    .X(_04958_));
 sky130_vsdinv _27246_ (.A(_04952_),
    .Y(_04959_));
 sky130_fd_sc_hd__or2_1 _27247_ (.A(_04959_),
    .B(_04954_),
    .X(_04960_));
 sky130_fd_sc_hd__or2_1 _27248_ (.A(_04958_),
    .B(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__nand2_1 _27249_ (.A(_04960_),
    .B(_04958_),
    .Y(_04962_));
 sky130_fd_sc_hd__and2_1 _27250_ (.A(_04961_),
    .B(_04962_),
    .X(_02598_));
 sky130_fd_sc_hd__or2_1 _27251_ (.A(_02366_),
    .B(_04956_),
    .X(_04963_));
 sky130_fd_sc_hd__nand2_1 _27252_ (.A(_04956_),
    .B(_02366_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand2_1 _27253_ (.A(_04963_),
    .B(_04964_),
    .Y(_02367_));
 sky130_fd_sc_hd__nor2_1 _27254_ (.A(_19800_),
    .B(_02368_),
    .Y(_04965_));
 sky130_fd_sc_hd__and2_1 _27255_ (.A(net314),
    .B(_02368_),
    .X(_04966_));
 sky130_fd_sc_hd__nor2_1 _27256_ (.A(_04965_),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__a21bo_1 _27257_ (.A1(_19801_),
    .A2(_02365_),
    .B1_N(_04962_),
    .X(_04968_));
 sky130_fd_sc_hd__xor2_1 _27258_ (.A(_04967_),
    .B(_04968_),
    .X(_02599_));
 sky130_fd_sc_hd__nor2_1 _27259_ (.A(net347),
    .B(_04964_),
    .Y(_04969_));
 sky130_fd_sc_hd__and2_1 _27260_ (.A(_04964_),
    .B(_19435_),
    .X(_04970_));
 sky130_fd_sc_hd__or2_1 _27261_ (.A(_04969_),
    .B(_04970_),
    .X(_02370_));
 sky130_fd_sc_hd__and2_1 _27262_ (.A(_04958_),
    .B(_04967_),
    .X(_04971_));
 sky130_fd_sc_hd__o21ai_1 _27263_ (.A1(_04959_),
    .A2(_04954_),
    .B1(_04971_),
    .Y(_04972_));
 sky130_vsdinv _27264_ (.A(_04965_),
    .Y(_04973_));
 sky130_fd_sc_hd__a31oi_2 _27265_ (.A1(_04973_),
    .A2(net313),
    .A3(_02365_),
    .B1(_04966_),
    .Y(_04974_));
 sky130_fd_sc_hd__or2_1 _27266_ (.A(net315),
    .B(_02371_),
    .X(_04975_));
 sky130_fd_sc_hd__nand2_1 _27267_ (.A(net315),
    .B(_02371_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2_1 _27268_ (.A(_04975_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__a21oi_2 _27269_ (.A1(_04972_),
    .A2(_04974_),
    .B1(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__and3_1 _27270_ (.A(_04972_),
    .B(_04977_),
    .C(_04974_),
    .X(_04979_));
 sky130_fd_sc_hd__nor2_1 _27271_ (.A(_04978_),
    .B(_04979_),
    .Y(_02600_));
 sky130_fd_sc_hd__or2_1 _27272_ (.A(_02372_),
    .B(_04969_),
    .X(_04980_));
 sky130_fd_sc_hd__nand2_1 _27273_ (.A(_04969_),
    .B(_02372_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand2_1 _27274_ (.A(_04980_),
    .B(_04981_),
    .Y(_02373_));
 sky130_vsdinv _27275_ (.A(_04976_),
    .Y(_04982_));
 sky130_fd_sc_hd__or2_1 _27276_ (.A(net316),
    .B(_02374_),
    .X(_04983_));
 sky130_fd_sc_hd__nand2_1 _27277_ (.A(net316),
    .B(_02374_),
    .Y(_04984_));
 sky130_fd_sc_hd__and2_1 _27278_ (.A(_04983_),
    .B(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__or3_2 _27279_ (.A(_04982_),
    .B(_04985_),
    .C(_04978_),
    .X(_04986_));
 sky130_fd_sc_hd__o21ai_2 _27280_ (.A1(_04982_),
    .A2(_04978_),
    .B1(_04985_),
    .Y(_04987_));
 sky130_fd_sc_hd__and2_1 _27281_ (.A(_04986_),
    .B(_04987_),
    .X(_02601_));
 sky130_fd_sc_hd__nor2_1 _27282_ (.A(net350),
    .B(_04981_),
    .Y(_04988_));
 sky130_vsdinv _27283_ (.A(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__nand2_1 _27284_ (.A(_04981_),
    .B(net350),
    .Y(_04990_));
 sky130_fd_sc_hd__nand2_1 _27285_ (.A(_04989_),
    .B(_04990_),
    .Y(_02376_));
 sky130_fd_sc_hd__or2_1 _27286_ (.A(net318),
    .B(_02377_),
    .X(_04991_));
 sky130_fd_sc_hd__nand2_1 _27287_ (.A(_19796_),
    .B(_02377_),
    .Y(_04992_));
 sky130_fd_sc_hd__nand2_1 _27288_ (.A(_04991_),
    .B(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__a21oi_2 _27289_ (.A1(_04987_),
    .A2(_04984_),
    .B1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__and3_1 _27290_ (.A(_04987_),
    .B(_04984_),
    .C(_04993_),
    .X(_04995_));
 sky130_fd_sc_hd__nor2_1 _27291_ (.A(_04994_),
    .B(_04995_),
    .Y(_02603_));
 sky130_fd_sc_hd__nand2_1 _27292_ (.A(_04989_),
    .B(_19433_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_1 _27293_ (.A(_04988_),
    .B(_02378_),
    .Y(_04997_));
 sky130_fd_sc_hd__nand2_1 _27294_ (.A(_04996_),
    .B(_04997_),
    .Y(_02379_));
 sky130_vsdinv _27295_ (.A(_04992_),
    .Y(_04998_));
 sky130_fd_sc_hd__or2_1 _27296_ (.A(net319),
    .B(_02380_),
    .X(_04999_));
 sky130_fd_sc_hd__nand2_2 _27297_ (.A(net319),
    .B(_02380_),
    .Y(_05000_));
 sky130_fd_sc_hd__and2_1 _27298_ (.A(_04999_),
    .B(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__or3_2 _27299_ (.A(_04998_),
    .B(_05001_),
    .C(_04994_),
    .X(_05002_));
 sky130_fd_sc_hd__o21ai_2 _27300_ (.A1(_04998_),
    .A2(_04994_),
    .B1(_05001_),
    .Y(_05003_));
 sky130_fd_sc_hd__and2_1 _27301_ (.A(_05002_),
    .B(_05003_),
    .X(_02604_));
 sky130_fd_sc_hd__or2_1 _27302_ (.A(_19432_),
    .B(_04997_),
    .X(_05004_));
 sky130_fd_sc_hd__nand2_1 _27303_ (.A(_04997_),
    .B(_19432_),
    .Y(_05005_));
 sky130_fd_sc_hd__nand2_1 _27304_ (.A(_05004_),
    .B(_05005_),
    .Y(_02382_));
 sky130_fd_sc_hd__or2_1 _27305_ (.A(net320),
    .B(_02383_),
    .X(_05006_));
 sky130_fd_sc_hd__nand2_1 _27306_ (.A(_19794_),
    .B(_02383_),
    .Y(_05007_));
 sky130_fd_sc_hd__nand2_2 _27307_ (.A(_05006_),
    .B(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__a21oi_4 _27308_ (.A1(_05003_),
    .A2(_05000_),
    .B1(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__and3_1 _27309_ (.A(_05003_),
    .B(_05000_),
    .C(_05008_),
    .X(_05010_));
 sky130_fd_sc_hd__nor2_1 _27310_ (.A(_05009_),
    .B(_05010_),
    .Y(_02605_));
 sky130_fd_sc_hd__nor2_1 _27311_ (.A(_19431_),
    .B(_05004_),
    .Y(_05011_));
 sky130_fd_sc_hd__and2_1 _27312_ (.A(_05004_),
    .B(_19431_),
    .X(_05012_));
 sky130_fd_sc_hd__or2_1 _27313_ (.A(_05011_),
    .B(_05012_),
    .X(_02385_));
 sky130_vsdinv _27314_ (.A(_05007_),
    .Y(_05013_));
 sky130_fd_sc_hd__or2_1 _27315_ (.A(net321),
    .B(_02386_),
    .X(_05014_));
 sky130_fd_sc_hd__nand2_1 _27316_ (.A(_19793_),
    .B(_02386_),
    .Y(_05015_));
 sky130_fd_sc_hd__and2_1 _27317_ (.A(_05014_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__or3_2 _27318_ (.A(_05013_),
    .B(_05016_),
    .C(_05009_),
    .X(_05017_));
 sky130_fd_sc_hd__o21ai_2 _27319_ (.A1(_05013_),
    .A2(_05009_),
    .B1(_05016_),
    .Y(_05018_));
 sky130_fd_sc_hd__and2_1 _27320_ (.A(_05017_),
    .B(_05018_),
    .X(_02606_));
 sky130_fd_sc_hd__or2_1 _27321_ (.A(_02387_),
    .B(_05011_),
    .X(_05019_));
 sky130_fd_sc_hd__nand2_1 _27322_ (.A(_05011_),
    .B(_02387_),
    .Y(_05020_));
 sky130_fd_sc_hd__nand2_1 _27323_ (.A(_05019_),
    .B(_05020_),
    .Y(_02388_));
 sky130_fd_sc_hd__or2_1 _27324_ (.A(_19792_),
    .B(_02389_),
    .X(_05021_));
 sky130_fd_sc_hd__nand2_1 _27325_ (.A(_19792_),
    .B(_02389_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand2_1 _27326_ (.A(_05021_),
    .B(_05022_),
    .Y(_05023_));
 sky130_vsdinv _27327_ (.A(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_1 _27328_ (.A(_05018_),
    .B(_05015_),
    .Y(_05025_));
 sky130_fd_sc_hd__or2_1 _27329_ (.A(_05024_),
    .B(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__nand2_1 _27330_ (.A(_05025_),
    .B(_05024_),
    .Y(_05027_));
 sky130_fd_sc_hd__and2_1 _27331_ (.A(_05026_),
    .B(_05027_),
    .X(_02607_));
 sky130_fd_sc_hd__nor2_1 _27332_ (.A(net355),
    .B(_05020_),
    .Y(_05028_));
 sky130_vsdinv _27333_ (.A(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__nand2_1 _27334_ (.A(_05020_),
    .B(net355),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2_1 _27335_ (.A(_05029_),
    .B(_05030_),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_1 _27336_ (.A(_19790_),
    .B(_02392_),
    .Y(_05031_));
 sky130_fd_sc_hd__nand2_1 _27337_ (.A(_19790_),
    .B(_02392_),
    .Y(_05032_));
 sky130_fd_sc_hd__or2b_1 _27338_ (.A(_05031_),
    .B_N(_05032_),
    .X(_05033_));
 sky130_vsdinv _27339_ (.A(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand2_1 _27340_ (.A(_05027_),
    .B(_05022_),
    .Y(_05035_));
 sky130_fd_sc_hd__xor2_1 _27341_ (.A(_05034_),
    .B(_05035_),
    .X(_02608_));
 sky130_fd_sc_hd__nand2_1 _27342_ (.A(_05029_),
    .B(net356),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_1 _27343_ (.A(_05028_),
    .B(_02393_),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2_1 _27344_ (.A(_05036_),
    .B(_05037_),
    .Y(_02394_));
 sky130_fd_sc_hd__nor2_1 _27345_ (.A(net324),
    .B(_02395_),
    .Y(_05038_));
 sky130_vsdinv _27346_ (.A(_02395_),
    .Y(_05039_));
 sky130_fd_sc_hd__nor2_1 _27347_ (.A(_20210_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__nor2_1 _27348_ (.A(_05038_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__nand2_1 _27349_ (.A(_05034_),
    .B(_05024_),
    .Y(_05042_));
 sky130_fd_sc_hd__a21oi_2 _27350_ (.A1(_05018_),
    .A2(_05015_),
    .B1(_05042_),
    .Y(_05043_));
 sky130_vsdinv _27351_ (.A(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__o21a_1 _27352_ (.A1(_05022_),
    .A2(_05031_),
    .B1(_05032_),
    .X(_05045_));
 sky130_fd_sc_hd__nand2_1 _27353_ (.A(_05044_),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__or2_1 _27354_ (.A(_05041_),
    .B(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__nand2_1 _27355_ (.A(_05046_),
    .B(_05041_),
    .Y(_05048_));
 sky130_fd_sc_hd__and2_1 _27356_ (.A(_05047_),
    .B(_05048_),
    .X(_02609_));
 sky130_fd_sc_hd__nor2_1 _27357_ (.A(_19429_),
    .B(_05037_),
    .Y(_05049_));
 sky130_fd_sc_hd__and2_1 _27358_ (.A(_05037_),
    .B(_19429_),
    .X(_05050_));
 sky130_fd_sc_hd__or2_1 _27359_ (.A(_05049_),
    .B(_05050_),
    .X(_02397_));
 sky130_fd_sc_hd__nor2_1 _27360_ (.A(_19789_),
    .B(_02398_),
    .Y(_05051_));
 sky130_vsdinv _27361_ (.A(_02398_),
    .Y(_05052_));
 sky130_fd_sc_hd__nor2_1 _27362_ (.A(_20655_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__nor2_2 _27363_ (.A(_05051_),
    .B(_05053_),
    .Y(_05054_));
 sky130_vsdinv _27364_ (.A(_05040_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_1 _27365_ (.A(_05048_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__xor2_1 _27366_ (.A(_05054_),
    .B(_05056_),
    .X(_02610_));
 sky130_fd_sc_hd__or2_1 _27367_ (.A(_02399_),
    .B(_05049_),
    .X(_05057_));
 sky130_fd_sc_hd__and4_2 _27368_ (.A(_05028_),
    .B(_02399_),
    .C(_02396_),
    .D(_02393_),
    .X(_05058_));
 sky130_vsdinv _27369_ (.A(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_1 _27370_ (.A(_05057_),
    .B(_05059_),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _27371_ (.A(net326),
    .B(_02401_),
    .Y(_05060_));
 sky130_vsdinv _27372_ (.A(_02401_),
    .Y(_05061_));
 sky130_fd_sc_hd__nor2_4 _27373_ (.A(_20236_),
    .B(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__nor2_1 _27374_ (.A(_05060_),
    .B(_05062_),
    .Y(_05063_));
 sky130_vsdinv _27375_ (.A(_05045_),
    .Y(_05064_));
 sky130_fd_sc_hd__nand2_1 _27376_ (.A(_05041_),
    .B(_05054_),
    .Y(_05065_));
 sky130_fd_sc_hd__o21bai_2 _27377_ (.A1(_05064_),
    .A2(_05043_),
    .B1_N(_05065_),
    .Y(_05066_));
 sky130_vsdinv _27378_ (.A(_05053_),
    .Y(_05067_));
 sky130_fd_sc_hd__o21a_1 _27379_ (.A1(_05051_),
    .A2(_05055_),
    .B1(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_1 _27380_ (.A(_05066_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__xor2_1 _27381_ (.A(_05063_),
    .B(_05069_),
    .X(_02611_));
 sky130_fd_sc_hd__nand2_1 _27382_ (.A(_05059_),
    .B(net359),
    .Y(_05070_));
 sky130_fd_sc_hd__nand2_1 _27383_ (.A(_05058_),
    .B(_02402_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _27384_ (.A(_05070_),
    .B(_05071_),
    .Y(_02403_));
 sky130_vsdinv _27385_ (.A(_02404_),
    .Y(_05072_));
 sky130_fd_sc_hd__nor2_1 _27386_ (.A(_20231_),
    .B(_05072_),
    .Y(_05073_));
 sky130_vsdinv _27387_ (.A(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand2_1 _27388_ (.A(_20231_),
    .B(_05072_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand2_1 _27389_ (.A(_05074_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__a22oi_4 _27390_ (.A1(_20236_),
    .A2(_05061_),
    .B1(_05066_),
    .B2(_05068_),
    .Y(_05077_));
 sky130_fd_sc_hd__or3_2 _27391_ (.A(_05062_),
    .B(_05076_),
    .C(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__o21ai_1 _27392_ (.A1(_05062_),
    .A2(_05077_),
    .B1(_05076_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand2_1 _27393_ (.A(_05078_),
    .B(_05079_),
    .Y(_02612_));
 sky130_fd_sc_hd__nand2_1 _27394_ (.A(_05071_),
    .B(_19428_),
    .Y(_05080_));
 sky130_fd_sc_hd__nor2_2 _27395_ (.A(_19428_),
    .B(net359),
    .Y(_05081_));
 sky130_fd_sc_hd__nand2_1 _27396_ (.A(_05058_),
    .B(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__nand2_1 _27397_ (.A(_05080_),
    .B(_05082_),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _27398_ (.A(_19787_),
    .B(_02407_),
    .Y(_05083_));
 sky130_vsdinv _27399_ (.A(_02407_),
    .Y(_05084_));
 sky130_fd_sc_hd__nor2_1 _27400_ (.A(_20678_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__nor2_1 _27401_ (.A(_05083_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__o22ai_4 _27402_ (.A1(_19788_),
    .A2(_02404_),
    .B1(_05062_),
    .B2(_05077_),
    .Y(_05087_));
 sky130_fd_sc_hd__nand2_1 _27403_ (.A(_05087_),
    .B(_05074_),
    .Y(_05088_));
 sky130_fd_sc_hd__xor2_1 _27404_ (.A(_05086_),
    .B(_05088_),
    .X(_02614_));
 sky130_fd_sc_hd__a21o_1 _27405_ (.A1(_05058_),
    .A2(_05081_),
    .B1(_18471_),
    .X(_05089_));
 sky130_fd_sc_hd__nand3_1 _27406_ (.A(_05058_),
    .B(_18471_),
    .C(_05081_),
    .Y(_05090_));
 sky130_fd_sc_hd__nand2_1 _27407_ (.A(_05089_),
    .B(_05090_),
    .Y(_02408_));
 sky130_fd_sc_hd__nor2_1 _27408_ (.A(_02409_),
    .B(_20684_),
    .Y(_05091_));
 sky130_fd_sc_hd__and2_1 _27409_ (.A(_20684_),
    .B(_02409_),
    .X(_05092_));
 sky130_fd_sc_hd__a22oi_1 _27410_ (.A1(_20678_),
    .A2(_05084_),
    .B1(_05087_),
    .B2(_05074_),
    .Y(_05093_));
 sky130_fd_sc_hd__o22ai_1 _27411_ (.A1(_05091_),
    .A2(_05092_),
    .B1(_05085_),
    .B2(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__nor2_1 _27412_ (.A(_05091_),
    .B(_05092_),
    .Y(_05095_));
 sky130_fd_sc_hd__o2bb2ai_1 _27413_ (.A1_N(_05074_),
    .A2_N(_05087_),
    .B1(_19787_),
    .B2(_02407_),
    .Y(_05096_));
 sky130_fd_sc_hd__o211ai_1 _27414_ (.A1(_20678_),
    .A2(_05084_),
    .B1(_05095_),
    .C1(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__nand2_1 _27415_ (.A(_05094_),
    .B(_05097_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _27416_ (.A(_19687_),
    .B(_19931_),
    .Y(_05098_));
 sky130_fd_sc_hd__nand2_1 _27417_ (.A(_19684_),
    .B(_19934_),
    .Y(_05099_));
 sky130_fd_sc_hd__nor2_4 _27418_ (.A(_05098_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__and2_2 _27419_ (.A(_05098_),
    .B(_05099_),
    .X(_05101_));
 sky130_fd_sc_hd__nor2_8 _27420_ (.A(_05100_),
    .B(_05101_),
    .Y(_02624_));
 sky130_vsdinv _27421_ (.A(_05100_),
    .Y(_05102_));
 sky130_fd_sc_hd__nand2_1 _27422_ (.A(_19687_),
    .B(_19928_),
    .Y(_05103_));
 sky130_fd_sc_hd__nand2_1 _27423_ (.A(_19680_),
    .B(_19684_),
    .Y(_05104_));
 sky130_fd_sc_hd__buf_4 _27424_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05105_));
 sky130_vsdinv _27425_ (.A(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__or3_1 _27426_ (.A(_05104_),
    .B(_05106_),
    .C(net453),
    .X(_05107_));
 sky130_fd_sc_hd__a22o_1 _27427_ (.A1(_19680_),
    .A2(_19934_),
    .B1(_19684_),
    .B2(_19931_),
    .X(_05108_));
 sky130_fd_sc_hd__nand2_1 _27428_ (.A(_05107_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__or2_1 _27429_ (.A(_05103_),
    .B(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__nand2_1 _27430_ (.A(_05109_),
    .B(_05103_),
    .Y(_05111_));
 sky130_fd_sc_hd__nand2_1 _27431_ (.A(_05110_),
    .B(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__nor2_2 _27432_ (.A(_05102_),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__and2_1 _27433_ (.A(_05112_),
    .B(_05102_),
    .X(_05114_));
 sky130_fd_sc_hd__nor2_1 _27434_ (.A(_05113_),
    .B(_05114_),
    .Y(_02625_));
 sky130_fd_sc_hd__o21a_1 _27435_ (.A1(_05103_),
    .A2(_05109_),
    .B1(_05107_),
    .X(_05115_));
 sky130_fd_sc_hd__clkbuf_4 _27436_ (.A(\pcpi_mul.rs2[2] ),
    .X(_05116_));
 sky130_fd_sc_hd__buf_4 _27437_ (.A(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__clkbuf_4 _27438_ (.A(\pcpi_mul.rs2[1] ),
    .X(_05118_));
 sky130_fd_sc_hd__buf_4 _27439_ (.A(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__buf_4 _27440_ (.A(_19926_),
    .X(_05120_));
 sky130_fd_sc_hd__buf_6 _27441_ (.A(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__buf_4 _27442_ (.A(\pcpi_mul.rs1[1] ),
    .X(_05122_));
 sky130_fd_sc_hd__buf_4 _27443_ (.A(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__and4_2 _27444_ (.A(_05117_),
    .B(_05119_),
    .C(_05121_),
    .D(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__clkbuf_4 _27445_ (.A(_19678_),
    .X(_05125_));
 sky130_fd_sc_hd__clkbuf_4 _27446_ (.A(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__buf_6 _27447_ (.A(_19926_),
    .X(_05127_));
 sky130_fd_sc_hd__buf_6 _27448_ (.A(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__a22o_2 _27449_ (.A1(_05126_),
    .A2(_05123_),
    .B1(_19683_),
    .B2(_05128_),
    .X(_05129_));
 sky130_vsdinv _27450_ (.A(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__buf_6 _27451_ (.A(\pcpi_mul.rs2[3] ),
    .X(_05131_));
 sky130_fd_sc_hd__clkinv_8 _27452_ (.A(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__nor2_8 _27453_ (.A(_05132_),
    .B(_04840_),
    .Y(_05133_));
 sky130_fd_sc_hd__o21bai_2 _27454_ (.A1(_05124_),
    .A2(_05130_),
    .B1_N(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand3b_4 _27455_ (.A_N(_05124_),
    .B(_05129_),
    .C(_05133_),
    .Y(_05135_));
 sky130_fd_sc_hd__nand2_1 _27456_ (.A(_19687_),
    .B(_19925_),
    .Y(_05136_));
 sky130_fd_sc_hd__a21bo_1 _27457_ (.A1(_05134_),
    .A2(_05135_),
    .B1_N(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__nand3b_4 _27458_ (.A_N(_05136_),
    .B(_05134_),
    .C(_05135_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_1 _27459_ (.A(_05137_),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__or2_1 _27460_ (.A(_05115_),
    .B(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__nand2_1 _27461_ (.A(_05139_),
    .B(_05115_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_1 _27462_ (.A(_05140_),
    .B(_05141_),
    .Y(_05142_));
 sky130_vsdinv _27463_ (.A(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__or2_1 _27464_ (.A(_05113_),
    .B(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__nand2_1 _27465_ (.A(_05143_),
    .B(_05113_),
    .Y(_05145_));
 sky130_fd_sc_hd__and2_1 _27466_ (.A(_05144_),
    .B(_05145_),
    .X(_02626_));
 sky130_fd_sc_hd__buf_4 _27467_ (.A(_19922_),
    .X(_05146_));
 sky130_fd_sc_hd__clkbuf_4 _27468_ (.A(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__and4_4 _27469_ (.A(_05126_),
    .B(_19683_),
    .C(_05147_),
    .D(_05128_),
    .X(_05148_));
 sky130_vsdinv _27470_ (.A(_05126_),
    .Y(_05149_));
 sky130_fd_sc_hd__clkinv_8 _27471_ (.A(_19926_),
    .Y(_05150_));
 sky130_fd_sc_hd__buf_6 _27472_ (.A(_05150_),
    .X(_05151_));
 sky130_fd_sc_hd__buf_6 _27473_ (.A(_19681_),
    .X(_05152_));
 sky130_vsdinv _27474_ (.A(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__inv_8 _27475_ (.A(_19922_),
    .Y(_05154_));
 sky130_fd_sc_hd__buf_6 _27476_ (.A(_05154_),
    .X(_05155_));
 sky130_fd_sc_hd__o22a_4 _27477_ (.A1(_05149_),
    .A2(_05151_),
    .B1(_05153_),
    .B2(_05155_),
    .X(_05156_));
 sky130_fd_sc_hd__buf_6 _27478_ (.A(_05131_),
    .X(_05157_));
 sky130_fd_sc_hd__buf_6 _27479_ (.A(_19930_),
    .X(_05158_));
 sky130_fd_sc_hd__nand2_4 _27480_ (.A(_05157_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__o21ai_4 _27481_ (.A1(_05148_),
    .A2(_05156_),
    .B1(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__buf_6 _27482_ (.A(_19678_),
    .X(_05161_));
 sky130_fd_sc_hd__buf_4 _27483_ (.A(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__buf_6 _27484_ (.A(_05118_),
    .X(_05163_));
 sky130_fd_sc_hd__buf_4 _27485_ (.A(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__a22o_2 _27486_ (.A1(_05162_),
    .A2(_19928_),
    .B1(_05164_),
    .B2(_19925_),
    .X(_05165_));
 sky130_vsdinv _27487_ (.A(_05159_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand3b_4 _27488_ (.A_N(_05148_),
    .B(_05165_),
    .C(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__clkbuf_4 _27489_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05168_));
 sky130_fd_sc_hd__clkbuf_4 _27490_ (.A(_05168_),
    .X(_05169_));
 sky130_fd_sc_hd__nand2_1 _27491_ (.A(_05169_),
    .B(_19933_),
    .Y(_05170_));
 sky130_fd_sc_hd__buf_6 _27492_ (.A(_19685_),
    .X(_05171_));
 sky130_fd_sc_hd__buf_4 _27493_ (.A(\pcpi_mul.rs1[4] ),
    .X(_05172_));
 sky130_fd_sc_hd__buf_4 _27494_ (.A(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__buf_6 _27495_ (.A(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__nand2_2 _27496_ (.A(_05171_),
    .B(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__nor2_2 _27497_ (.A(_05170_),
    .B(_05175_),
    .Y(_05176_));
 sky130_vsdinv _27498_ (.A(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__nand2_1 _27499_ (.A(_05170_),
    .B(_05175_),
    .Y(_05178_));
 sky130_fd_sc_hd__and2_2 _27500_ (.A(_05177_),
    .B(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__a21oi_4 _27501_ (.A1(_05160_),
    .A2(_05167_),
    .B1(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__nand2_1 _27502_ (.A(_05177_),
    .B(_05178_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _27503_ (.A(_05160_),
    .B(_05167_),
    .Y(_05182_));
 sky130_fd_sc_hd__nor2_2 _27504_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__o21ai_4 _27505_ (.A1(_05180_),
    .A2(_05183_),
    .B1(_05138_),
    .Y(_05184_));
 sky130_fd_sc_hd__nand2_1 _27506_ (.A(_05182_),
    .B(_05181_),
    .Y(_05185_));
 sky130_fd_sc_hd__nand3_4 _27507_ (.A(_05179_),
    .B(_05167_),
    .C(_05160_),
    .Y(_05186_));
 sky130_fd_sc_hd__nand3b_4 _27508_ (.A_N(_05138_),
    .B(_05185_),
    .C(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__a21oi_2 _27509_ (.A1(_05133_),
    .A2(_05129_),
    .B1(_05124_),
    .Y(_05188_));
 sky130_vsdinv _27510_ (.A(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__a21o_1 _27511_ (.A1(_05184_),
    .A2(_05187_),
    .B1(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__nand3_2 _27512_ (.A(_05184_),
    .B(_05189_),
    .C(_05187_),
    .Y(_05191_));
 sky130_fd_sc_hd__nand2_1 _27513_ (.A(_05190_),
    .B(_05191_),
    .Y(_05192_));
 sky130_vsdinv _27514_ (.A(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__nand2_1 _27515_ (.A(_05145_),
    .B(_05140_),
    .Y(_05194_));
 sky130_fd_sc_hd__or2_1 _27516_ (.A(_05193_),
    .B(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__nand2_1 _27517_ (.A(_05194_),
    .B(_05193_),
    .Y(_05196_));
 sky130_fd_sc_hd__and2_1 _27518_ (.A(_05195_),
    .B(_05196_),
    .X(_02627_));
 sky130_fd_sc_hd__buf_8 _27519_ (.A(_19669_),
    .X(_05197_));
 sky130_fd_sc_hd__clkbuf_8 _27520_ (.A(\pcpi_mul.rs1[0] ),
    .X(_05198_));
 sky130_fd_sc_hd__buf_6 _27521_ (.A(_19929_),
    .X(_05199_));
 sky130_fd_sc_hd__a22oi_4 _27522_ (.A1(_05197_),
    .A2(_05198_),
    .B1(_05169_),
    .B2(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__buf_6 _27523_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05201_));
 sky130_fd_sc_hd__nand2_2 _27524_ (.A(_05201_),
    .B(_05105_),
    .Y(_05202_));
 sky130_fd_sc_hd__buf_6 _27525_ (.A(_19669_),
    .X(_05203_));
 sky130_fd_sc_hd__clkbuf_4 _27526_ (.A(\pcpi_mul.rs1[0] ),
    .X(_05204_));
 sky130_fd_sc_hd__nand2_2 _27527_ (.A(_05203_),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__nor2_4 _27528_ (.A(_05202_),
    .B(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__buf_1 _27529_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05207_));
 sky130_fd_sc_hd__clkbuf_8 _27530_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05208_));
 sky130_fd_sc_hd__nand2_4 _27531_ (.A(_05207_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__o21ai_2 _27532_ (.A1(_05200_),
    .A2(_05206_),
    .B1(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__buf_6 _27533_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05211_));
 sky130_fd_sc_hd__clkbuf_4 _27534_ (.A(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__buf_8 _27535_ (.A(_19932_),
    .X(_05213_));
 sky130_fd_sc_hd__nand3b_4 _27536_ (.A_N(_05202_),
    .B(_05212_),
    .C(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__nand2_2 _27537_ (.A(_05202_),
    .B(_05205_),
    .Y(_05215_));
 sky130_vsdinv _27538_ (.A(_05209_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand3_2 _27539_ (.A(_05214_),
    .B(_05215_),
    .C(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__nand3_4 _27540_ (.A(_05210_),
    .B(_05217_),
    .C(_05176_),
    .Y(_05218_));
 sky130_fd_sc_hd__o21ai_2 _27541_ (.A1(_05200_),
    .A2(_05206_),
    .B1(_05216_),
    .Y(_05219_));
 sky130_fd_sc_hd__nand3_2 _27542_ (.A(_05214_),
    .B(_05215_),
    .C(_05209_),
    .Y(_05220_));
 sky130_fd_sc_hd__nand3_4 _27543_ (.A(_05219_),
    .B(_05220_),
    .C(_05177_),
    .Y(_05221_));
 sky130_fd_sc_hd__nand2_1 _27544_ (.A(_05218_),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__clkbuf_8 _27545_ (.A(_05152_),
    .X(_05223_));
 sky130_fd_sc_hd__buf_6 _27546_ (.A(_05172_),
    .X(_05224_));
 sky130_fd_sc_hd__buf_6 _27547_ (.A(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__a22oi_4 _27548_ (.A1(_05126_),
    .A2(_05147_),
    .B1(_05223_),
    .B2(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__buf_6 _27549_ (.A(_05118_),
    .X(_05227_));
 sky130_fd_sc_hd__and4_4 _27550_ (.A(_19679_),
    .B(_05227_),
    .C(_05174_),
    .D(_19924_),
    .X(_05228_));
 sky130_fd_sc_hd__buf_6 _27551_ (.A(\pcpi_mul.rs1[2] ),
    .X(_05229_));
 sky130_fd_sc_hd__buf_6 _27552_ (.A(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__nand2_4 _27553_ (.A(_19676_),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__o21bai_1 _27554_ (.A1(_05226_),
    .A2(_05228_),
    .B1_N(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__buf_6 _27555_ (.A(_05116_),
    .X(_05233_));
 sky130_fd_sc_hd__nand2_1 _27556_ (.A(_05233_),
    .B(_19924_),
    .Y(_05234_));
 sky130_fd_sc_hd__buf_6 _27557_ (.A(_19682_),
    .X(_05235_));
 sky130_fd_sc_hd__buf_4 _27558_ (.A(_19919_),
    .X(_05236_));
 sky130_fd_sc_hd__buf_6 _27559_ (.A(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__nand3b_4 _27560_ (.A_N(_05234_),
    .B(_05235_),
    .C(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__buf_4 _27561_ (.A(_19682_),
    .X(_05239_));
 sky130_fd_sc_hd__a22o_2 _27562_ (.A1(_05117_),
    .A2(_05147_),
    .B1(_05239_),
    .B2(_05225_),
    .X(_05240_));
 sky130_fd_sc_hd__nand3_1 _27563_ (.A(_05238_),
    .B(_05231_),
    .C(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__nand2_2 _27564_ (.A(_05232_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__nand2_2 _27565_ (.A(_05222_),
    .B(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__nand3b_4 _27566_ (.A_N(_05242_),
    .B(_05218_),
    .C(_05221_),
    .Y(_05244_));
 sky130_fd_sc_hd__a21o_1 _27567_ (.A1(_05243_),
    .A2(_05244_),
    .B1(_05186_),
    .X(_05245_));
 sky130_fd_sc_hd__nand3_4 _27568_ (.A(_05243_),
    .B(_05186_),
    .C(_05244_),
    .Y(_05246_));
 sky130_fd_sc_hd__nand2_1 _27569_ (.A(_05245_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__nor3_4 _27570_ (.A(_05148_),
    .B(_05159_),
    .C(_05156_),
    .Y(_05248_));
 sky130_fd_sc_hd__nor2_4 _27571_ (.A(_05148_),
    .B(_05248_),
    .Y(_05249_));
 sky130_vsdinv _27572_ (.A(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__nand2_2 _27573_ (.A(_05247_),
    .B(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand3_4 _27574_ (.A(_05245_),
    .B(_05246_),
    .C(_05249_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand2_1 _27575_ (.A(_05187_),
    .B(_05188_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2_2 _27576_ (.A(_05253_),
    .B(_05184_),
    .Y(_05254_));
 sky130_fd_sc_hd__a21oi_2 _27577_ (.A1(_05251_),
    .A2(_05252_),
    .B1(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__nor2_1 _27578_ (.A(_05115_),
    .B(_05139_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand3_2 _27579_ (.A(_05190_),
    .B(_05191_),
    .C(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__a31oi_2 _27580_ (.A1(_05254_),
    .A2(_05251_),
    .A3(_05252_),
    .B1(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__buf_4 _27581_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05259_));
 sky130_vsdinv _27582_ (.A(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__buf_8 _27583_ (.A(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__nand2_2 _27584_ (.A(_05238_),
    .B(_05231_),
    .Y(_05262_));
 sky130_fd_sc_hd__buf_6 _27585_ (.A(\pcpi_mul.rs1[3] ),
    .X(_05263_));
 sky130_fd_sc_hd__buf_6 _27586_ (.A(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_4 _27587_ (.A(_05131_),
    .B(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__buf_6 _27588_ (.A(_19678_),
    .X(_05266_));
 sky130_fd_sc_hd__buf_6 _27589_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05267_));
 sky130_fd_sc_hd__buf_6 _27590_ (.A(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__a22oi_4 _27591_ (.A1(_05266_),
    .A2(_05236_),
    .B1(_05152_),
    .B2(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__clkbuf_4 _27592_ (.A(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__buf_4 _27593_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05271_));
 sky130_fd_sc_hd__buf_6 _27594_ (.A(_05172_),
    .X(_05272_));
 sky130_fd_sc_hd__and4_1 _27595_ (.A(_05116_),
    .B(_05118_),
    .C(_05271_),
    .D(_05272_),
    .X(_05273_));
 sky130_fd_sc_hd__buf_2 _27596_ (.A(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__nor3_4 _27597_ (.A(_05265_),
    .B(_05270_),
    .C(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__o21a_1 _27598_ (.A1(_05270_),
    .A2(_05274_),
    .B1(_05265_),
    .X(_05276_));
 sky130_fd_sc_hd__buf_6 _27599_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05277_));
 sky130_fd_sc_hd__inv_4 _27600_ (.A(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__buf_2 _27601_ (.A(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__clkbuf_8 _27602_ (.A(_19669_),
    .X(_05280_));
 sky130_fd_sc_hd__buf_6 _27603_ (.A(_19929_),
    .X(_05281_));
 sky130_fd_sc_hd__buf_6 _27604_ (.A(_05168_),
    .X(_05282_));
 sky130_fd_sc_hd__a22oi_4 _27605_ (.A1(_05280_),
    .A2(_05281_),
    .B1(_05282_),
    .B2(_19927_),
    .Y(_05283_));
 sky130_fd_sc_hd__buf_6 _27606_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05284_));
 sky130_fd_sc_hd__buf_8 _27607_ (.A(\pcpi_mul.rs2[4] ),
    .X(_05285_));
 sky130_fd_sc_hd__nand3_4 _27608_ (.A(_05284_),
    .B(_05285_),
    .C(_05281_),
    .Y(_05286_));
 sky130_fd_sc_hd__nor2_4 _27609_ (.A(_05150_),
    .B(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__o22ai_4 _27610_ (.A1(net474),
    .A2(net452),
    .B1(_05283_),
    .B2(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__o21ai_2 _27611_ (.A1(_05209_),
    .A2(_05200_),
    .B1(_05214_),
    .Y(_05289_));
 sky130_fd_sc_hd__buf_8 _27612_ (.A(\pcpi_mul.rs2[0] ),
    .X(_05290_));
 sky130_fd_sc_hd__buf_6 _27613_ (.A(_19912_),
    .X(_05291_));
 sky130_fd_sc_hd__nand2_4 _27614_ (.A(_05290_),
    .B(_05291_),
    .Y(_05292_));
 sky130_vsdinv _27615_ (.A(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__buf_4 _27616_ (.A(\pcpi_mul.rs2[5] ),
    .X(_05294_));
 sky130_fd_sc_hd__buf_6 _27617_ (.A(_05294_),
    .X(_05295_));
 sky130_fd_sc_hd__a22o_1 _27618_ (.A1(_05295_),
    .A2(_05199_),
    .B1(_05169_),
    .B2(_05230_),
    .X(_05296_));
 sky130_fd_sc_hd__o211ai_2 _27619_ (.A1(_05151_),
    .A2(_05286_),
    .B1(_05293_),
    .C1(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand3_4 _27620_ (.A(_05288_),
    .B(_05289_),
    .C(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__o21ai_2 _27621_ (.A1(_05283_),
    .A2(_05287_),
    .B1(_05293_),
    .Y(_05299_));
 sky130_fd_sc_hd__a21oi_2 _27622_ (.A1(_05216_),
    .A2(_05215_),
    .B1(_05206_),
    .Y(_05300_));
 sky130_fd_sc_hd__o211ai_4 _27623_ (.A1(_05151_),
    .A2(_05286_),
    .B1(_05292_),
    .C1(_05296_),
    .Y(_05301_));
 sky130_fd_sc_hd__nand3_4 _27624_ (.A(_05299_),
    .B(_05300_),
    .C(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__a2bb2oi_2 _27625_ (.A1_N(_05275_),
    .A2_N(_05276_),
    .B1(_05298_),
    .B2(_05302_),
    .Y(_05303_));
 sky130_vsdinv _27626_ (.A(_05265_),
    .Y(_05304_));
 sky130_fd_sc_hd__nor3_2 _27627_ (.A(_05304_),
    .B(_05270_),
    .C(_05274_),
    .Y(_05305_));
 sky130_fd_sc_hd__o21a_1 _27628_ (.A1(_05270_),
    .A2(_05274_),
    .B1(_05304_),
    .X(_05306_));
 sky130_fd_sc_hd__o211a_1 _27629_ (.A1(_05305_),
    .A2(_05306_),
    .B1(_05298_),
    .C1(_05302_),
    .X(_05307_));
 sky130_fd_sc_hd__a21boi_2 _27630_ (.A1(_05221_),
    .A2(_05242_),
    .B1_N(_05218_),
    .Y(_05308_));
 sky130_fd_sc_hd__o21ai_4 _27631_ (.A1(_05303_),
    .A2(_05307_),
    .B1(_05308_),
    .Y(_05309_));
 sky130_vsdinv _27632_ (.A(_05269_),
    .Y(_05310_));
 sky130_fd_sc_hd__nand3b_1 _27633_ (.A_N(_05273_),
    .B(_05310_),
    .C(_05265_),
    .Y(_05311_));
 sky130_fd_sc_hd__o21ai_1 _27634_ (.A1(_05269_),
    .A2(_05274_),
    .B1(_05304_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand2_1 _27635_ (.A(_05311_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__a21o_1 _27636_ (.A1(_05302_),
    .A2(_05298_),
    .B1(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__nand2_1 _27637_ (.A(_05221_),
    .B(_05242_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand2_1 _27638_ (.A(_05315_),
    .B(_05218_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand3_2 _27639_ (.A(_05313_),
    .B(_05302_),
    .C(_05298_),
    .Y(_05317_));
 sky130_fd_sc_hd__nand3_4 _27640_ (.A(_05314_),
    .B(_05316_),
    .C(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__a22oi_4 _27641_ (.A1(_05240_),
    .A2(_05262_),
    .B1(_05309_),
    .B2(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__nor2_4 _27642_ (.A(_05231_),
    .B(_05226_),
    .Y(_05320_));
 sky130_fd_sc_hd__o211a_1 _27643_ (.A1(_05228_),
    .A2(_05320_),
    .B1(_05318_),
    .C1(_05309_),
    .X(_05321_));
 sky130_fd_sc_hd__o22ai_4 _27644_ (.A1(_05261_),
    .A2(_04842_),
    .B1(_05319_),
    .B2(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__nand2_2 _27645_ (.A(_05309_),
    .B(_05318_),
    .Y(_05323_));
 sky130_fd_sc_hd__nor2_8 _27646_ (.A(_05228_),
    .B(_05320_),
    .Y(_05324_));
 sky130_fd_sc_hd__nand2_2 _27647_ (.A(_05323_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand3b_4 _27648_ (.A_N(_05324_),
    .B(_05309_),
    .C(_05318_),
    .Y(_05326_));
 sky130_fd_sc_hd__nor2_4 _27649_ (.A(_05261_),
    .B(net453),
    .Y(_05327_));
 sky130_fd_sc_hd__nand3_4 _27650_ (.A(_05325_),
    .B(_05326_),
    .C(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hd__a21oi_1 _27651_ (.A1(_05243_),
    .A2(_05244_),
    .B1(_05186_),
    .Y(_05329_));
 sky130_fd_sc_hd__and2_1 _27652_ (.A(_05246_),
    .B(_05250_),
    .X(_05330_));
 sky130_fd_sc_hd__or2_2 _27653_ (.A(_05329_),
    .B(_05330_),
    .X(_05331_));
 sky130_fd_sc_hd__a21oi_2 _27654_ (.A1(_05322_),
    .A2(_05328_),
    .B1(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__o211a_1 _27655_ (.A1(_05329_),
    .A2(_05330_),
    .B1(_05328_),
    .C1(_05322_),
    .X(_05333_));
 sky130_fd_sc_hd__o22ai_2 _27656_ (.A1(_05255_),
    .A2(_05258_),
    .B1(_05332_),
    .B2(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__a21o_1 _27657_ (.A1(_05322_),
    .A2(_05328_),
    .B1(_05331_),
    .X(_05335_));
 sky130_fd_sc_hd__a21oi_2 _27658_ (.A1(_05247_),
    .A2(_05249_),
    .B1(_05254_),
    .Y(_05336_));
 sky130_fd_sc_hd__nand2_1 _27659_ (.A(_05330_),
    .B(_05245_),
    .Y(_05337_));
 sky130_fd_sc_hd__nand3_2 _27660_ (.A(_05251_),
    .B(_05254_),
    .C(_05252_),
    .Y(_05338_));
 sky130_fd_sc_hd__nor2_1 _27661_ (.A(_05181_),
    .B(_05248_),
    .Y(_05339_));
 sky130_fd_sc_hd__a21oi_2 _27662_ (.A1(_05339_),
    .A2(_05160_),
    .B1(_05180_),
    .Y(_05340_));
 sky130_vsdinv _27663_ (.A(_05115_),
    .Y(_05341_));
 sky130_fd_sc_hd__o2111ai_4 _27664_ (.A1(_05189_),
    .A2(_05340_),
    .B1(_05138_),
    .C1(_05137_),
    .D1(_05341_),
    .Y(_05342_));
 sky130_fd_sc_hd__a31oi_2 _27665_ (.A1(_05189_),
    .A2(_05187_),
    .A3(_05184_),
    .B1(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__a22oi_2 _27666_ (.A1(_05336_),
    .A2(_05337_),
    .B1(_05338_),
    .B2(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand3_4 _27667_ (.A(_05331_),
    .B(_05322_),
    .C(_05328_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand3_2 _27668_ (.A(_05335_),
    .B(_05344_),
    .C(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__nor2_1 _27669_ (.A(_05192_),
    .B(_05145_),
    .Y(_05347_));
 sky130_fd_sc_hd__nand2_1 _27670_ (.A(_05336_),
    .B(_05337_),
    .Y(_05348_));
 sky130_fd_sc_hd__and2_1 _27671_ (.A(_05348_),
    .B(_05338_),
    .X(_05349_));
 sky130_fd_sc_hd__nand2_1 _27672_ (.A(_05347_),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__a21oi_2 _27673_ (.A1(_05334_),
    .A2(_05346_),
    .B1(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__and3_1 _27674_ (.A(_05350_),
    .B(_05334_),
    .C(_05346_),
    .X(_05352_));
 sky130_fd_sc_hd__nor2_1 _27675_ (.A(_05351_),
    .B(_05352_),
    .Y(_02683_));
 sky130_fd_sc_hd__and3_1 _27676_ (.A(_05335_),
    .B(_05345_),
    .C(_05258_),
    .X(_05353_));
 sky130_fd_sc_hd__nor2_2 _27677_ (.A(_05348_),
    .B(_05332_),
    .Y(_05354_));
 sky130_fd_sc_hd__nand2_1 _27678_ (.A(_05313_),
    .B(_05302_),
    .Y(_05355_));
 sky130_fd_sc_hd__nand2_1 _27679_ (.A(_05355_),
    .B(_05298_),
    .Y(_05356_));
 sky130_fd_sc_hd__o22ai_4 _27680_ (.A1(_05151_),
    .A2(_05286_),
    .B1(_05292_),
    .B2(_05283_),
    .Y(_05357_));
 sky130_fd_sc_hd__clkbuf_8 _27681_ (.A(_05168_),
    .X(_05358_));
 sky130_fd_sc_hd__buf_6 _27682_ (.A(_05263_),
    .X(_05359_));
 sky130_fd_sc_hd__a22oi_4 _27683_ (.A1(_05280_),
    .A2(_05127_),
    .B1(_05358_),
    .B2(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__nand3_4 _27684_ (.A(_19669_),
    .B(_05168_),
    .C(_05229_),
    .Y(_05361_));
 sky130_fd_sc_hd__nor2_8 _27685_ (.A(_05154_),
    .B(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand2_4 _27686_ (.A(\pcpi_mul.rs2[0] ),
    .B(_19909_),
    .Y(_05363_));
 sky130_vsdinv _27687_ (.A(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__o21ai_2 _27688_ (.A1(_05360_),
    .A2(_05362_),
    .B1(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__buf_6 _27689_ (.A(_05168_),
    .X(_05366_));
 sky130_fd_sc_hd__a22o_2 _27690_ (.A1(_05284_),
    .A2(_05120_),
    .B1(_05366_),
    .B2(_05146_),
    .X(_05367_));
 sky130_fd_sc_hd__o211ai_4 _27691_ (.A1(_05155_),
    .A2(_05361_),
    .B1(_05363_),
    .C1(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__nand3b_4 _27692_ (.A_N(_05357_),
    .B(_05365_),
    .C(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__o21ai_4 _27693_ (.A1(_05360_),
    .A2(_05362_),
    .B1(_05363_),
    .Y(_05370_));
 sky130_fd_sc_hd__o211ai_4 _27694_ (.A1(_05154_),
    .A2(_05361_),
    .B1(_05364_),
    .C1(_05367_),
    .Y(_05371_));
 sky130_fd_sc_hd__nand3_4 _27695_ (.A(_05370_),
    .B(_05371_),
    .C(_05357_),
    .Y(_05372_));
 sky130_fd_sc_hd__nand2_1 _27696_ (.A(_05369_),
    .B(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hd__buf_8 _27697_ (.A(_05173_),
    .X(_05374_));
 sky130_fd_sc_hd__nand2_2 _27698_ (.A(_05131_),
    .B(_05374_),
    .Y(_05375_));
 sky130_vsdinv _27699_ (.A(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__buf_4 _27700_ (.A(\pcpi_mul.rs1[5] ),
    .X(_05377_));
 sky130_fd_sc_hd__buf_6 _27701_ (.A(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__buf_6 _27702_ (.A(\pcpi_mul.rs1[6] ),
    .X(_05379_));
 sky130_fd_sc_hd__buf_8 _27703_ (.A(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__a22oi_4 _27704_ (.A1(_05233_),
    .A2(_05378_),
    .B1(_05227_),
    .B2(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__buf_6 _27705_ (.A(_19681_),
    .X(_05382_));
 sky130_fd_sc_hd__clkbuf_8 _27706_ (.A(_05377_),
    .X(_05383_));
 sky130_fd_sc_hd__and4_4 _27707_ (.A(_05233_),
    .B(_05382_),
    .C(_05380_),
    .D(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__nor3_4 _27708_ (.A(_05376_),
    .B(_05381_),
    .C(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__o21a_1 _27709_ (.A1(_05381_),
    .A2(_05384_),
    .B1(_05376_),
    .X(_05386_));
 sky130_fd_sc_hd__nor2_4 _27710_ (.A(_05385_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__nand2_1 _27711_ (.A(_05373_),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__nor3_4 _27712_ (.A(_05375_),
    .B(_05381_),
    .C(_05384_),
    .Y(_05389_));
 sky130_fd_sc_hd__o21a_1 _27713_ (.A1(_05381_),
    .A2(_05384_),
    .B1(_05375_),
    .X(_05390_));
 sky130_fd_sc_hd__nor2_1 _27714_ (.A(_05389_),
    .B(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand3_2 _27715_ (.A(_05391_),
    .B(_05372_),
    .C(_05369_),
    .Y(_05392_));
 sky130_fd_sc_hd__nand3_4 _27716_ (.A(_05356_),
    .B(_05388_),
    .C(_05392_),
    .Y(_05393_));
 sky130_vsdinv _27717_ (.A(_05302_),
    .Y(_05394_));
 sky130_fd_sc_hd__o21a_1 _27718_ (.A1(_05275_),
    .A2(_05276_),
    .B1(_05298_),
    .X(_05395_));
 sky130_fd_sc_hd__a2bb2oi_4 _27719_ (.A1_N(_05389_),
    .A2_N(_05390_),
    .B1(_05372_),
    .B2(_05369_),
    .Y(_05396_));
 sky130_fd_sc_hd__o211a_1 _27720_ (.A1(_05385_),
    .A2(_05386_),
    .B1(_05372_),
    .C1(_05369_),
    .X(_05397_));
 sky130_fd_sc_hd__o22ai_4 _27721_ (.A1(_05394_),
    .A2(_05395_),
    .B1(_05396_),
    .B2(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__nor2_2 _27722_ (.A(_05304_),
    .B(_05274_),
    .Y(_05399_));
 sky130_fd_sc_hd__o2bb2ai_2 _27723_ (.A1_N(_05393_),
    .A2_N(_05398_),
    .B1(_05270_),
    .B2(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__nor2_2 _27724_ (.A(_05270_),
    .B(_05399_),
    .Y(_05401_));
 sky130_fd_sc_hd__nand3_2 _27725_ (.A(_05398_),
    .B(_05393_),
    .C(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__buf_2 _27726_ (.A(\pcpi_mul.rs2[7] ),
    .X(_05403_));
 sky130_fd_sc_hd__buf_4 _27727_ (.A(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__buf_6 _27728_ (.A(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__buf_6 _27729_ (.A(_05198_),
    .X(_05406_));
 sky130_fd_sc_hd__nand2_2 _27730_ (.A(_05405_),
    .B(_05406_),
    .Y(_05407_));
 sky130_fd_sc_hd__nand2_2 _27731_ (.A(_19668_),
    .B(_05158_),
    .Y(_05408_));
 sky130_fd_sc_hd__nor2_4 _27732_ (.A(_05407_),
    .B(_05408_),
    .Y(_05409_));
 sky130_vsdinv _27733_ (.A(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand2_1 _27734_ (.A(_05407_),
    .B(_05408_),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_2 _27735_ (.A(_05410_),
    .B(_05411_),
    .Y(_05412_));
 sky130_vsdinv _27736_ (.A(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__nand3_4 _27737_ (.A(_05400_),
    .B(_05402_),
    .C(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__nand2_1 _27738_ (.A(_05398_),
    .B(_05393_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand2_1 _27739_ (.A(_05415_),
    .B(_05401_),
    .Y(_05416_));
 sky130_fd_sc_hd__nand3b_2 _27740_ (.A_N(_05401_),
    .B(_05398_),
    .C(_05393_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand3_4 _27741_ (.A(_05416_),
    .B(_05412_),
    .C(_05417_),
    .Y(_05418_));
 sky130_vsdinv _27742_ (.A(_05327_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2_1 _27743_ (.A(_05325_),
    .B(_05326_),
    .Y(_05420_));
 sky130_fd_sc_hd__o2bb2ai_4 _27744_ (.A1_N(_05414_),
    .A2_N(_05418_),
    .B1(_05419_),
    .B2(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21oi_2 _27745_ (.A1(_05323_),
    .A2(_05324_),
    .B1(_05419_),
    .Y(_05422_));
 sky130_fd_sc_hd__o2111ai_4 _27746_ (.A1(_05324_),
    .A2(_05323_),
    .B1(_05422_),
    .C1(_05414_),
    .D1(_05418_),
    .Y(_05423_));
 sky130_fd_sc_hd__buf_2 _27747_ (.A(_05423_),
    .X(_05424_));
 sky130_vsdinv _27748_ (.A(_05318_),
    .Y(_05425_));
 sky130_fd_sc_hd__and3_1 _27749_ (.A(_05309_),
    .B(_05240_),
    .C(_05262_),
    .X(_05426_));
 sky130_fd_sc_hd__or2_2 _27750_ (.A(_05425_),
    .B(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__a21oi_2 _27751_ (.A1(_05421_),
    .A2(_05424_),
    .B1(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__o211a_1 _27752_ (.A1(_05425_),
    .A2(_05426_),
    .B1(_05424_),
    .C1(_05421_),
    .X(_05429_));
 sky130_fd_sc_hd__o22ai_2 _27753_ (.A1(_05333_),
    .A2(_05354_),
    .B1(_05428_),
    .B2(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__a21oi_1 _27754_ (.A1(_05335_),
    .A2(_05255_),
    .B1(_05333_),
    .Y(_05431_));
 sky130_fd_sc_hd__a21o_1 _27755_ (.A1(_05421_),
    .A2(_05424_),
    .B1(_05427_),
    .X(_05432_));
 sky130_fd_sc_hd__nand3_4 _27756_ (.A(_05421_),
    .B(_05424_),
    .C(_05427_),
    .Y(_05433_));
 sky130_fd_sc_hd__nand3_2 _27757_ (.A(_05431_),
    .B(_05432_),
    .C(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__nand2_1 _27758_ (.A(_05430_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__nor3_1 _27759_ (.A(_05351_),
    .B(_05353_),
    .C(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__o2bb2ai_1 _27760_ (.A1_N(_05434_),
    .A2_N(_05430_),
    .B1(_05353_),
    .B2(_05351_),
    .Y(_05437_));
 sky130_fd_sc_hd__nor2b_1 _27761_ (.A(_05436_),
    .B_N(_05437_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21oi_1 _27762_ (.A1(_05345_),
    .A2(_05433_),
    .B1(_05428_),
    .Y(_05438_));
 sky130_fd_sc_hd__buf_2 _27763_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05439_));
 sky130_fd_sc_hd__buf_6 _27764_ (.A(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__buf_4 _27765_ (.A(_19929_),
    .X(_05441_));
 sky130_fd_sc_hd__and4_4 _27766_ (.A(_05440_),
    .B(_19664_),
    .C(_05441_),
    .D(_05204_),
    .X(_05442_));
 sky130_fd_sc_hd__buf_6 _27767_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05443_));
 sky130_fd_sc_hd__nand2_2 _27768_ (.A(_05443_),
    .B(_05127_),
    .Y(_05444_));
 sky130_vsdinv _27769_ (.A(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__buf_4 _27770_ (.A(_05439_),
    .X(_05446_));
 sky130_fd_sc_hd__buf_6 _27771_ (.A(_05403_),
    .X(_05447_));
 sky130_fd_sc_hd__a22o_2 _27772_ (.A1(_05446_),
    .A2(_05204_),
    .B1(_05447_),
    .B2(_19930_),
    .X(_05448_));
 sky130_fd_sc_hd__nand3b_4 _27773_ (.A_N(_05442_),
    .B(_05445_),
    .C(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__buf_4 _27774_ (.A(\pcpi_mul.rs2[8] ),
    .X(_05450_));
 sky130_fd_sc_hd__buf_6 _27775_ (.A(_05450_),
    .X(_05451_));
 sky130_fd_sc_hd__buf_6 _27776_ (.A(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__a22oi_4 _27777_ (.A1(_05452_),
    .A2(_05406_),
    .B1(_05405_),
    .B2(_05158_),
    .Y(_05453_));
 sky130_fd_sc_hd__o21ai_4 _27778_ (.A1(_05453_),
    .A2(_05442_),
    .B1(_05444_),
    .Y(_05454_));
 sky130_fd_sc_hd__a21o_1 _27779_ (.A1(_05449_),
    .A2(_05454_),
    .B1(_05409_),
    .X(_05455_));
 sky130_fd_sc_hd__nand3_4 _27780_ (.A(_05449_),
    .B(_05409_),
    .C(_05454_),
    .Y(_05456_));
 sky130_fd_sc_hd__nand2_4 _27781_ (.A(_05455_),
    .B(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__a21oi_4 _27782_ (.A1(_05370_),
    .A2(_05371_),
    .B1(_05357_),
    .Y(_05458_));
 sky130_fd_sc_hd__o21ai_2 _27783_ (.A1(_05458_),
    .A2(_05387_),
    .B1(_05372_),
    .Y(_05459_));
 sky130_fd_sc_hd__nor2_2 _27784_ (.A(_05363_),
    .B(_05360_),
    .Y(_05460_));
 sky130_fd_sc_hd__nand2_2 _27785_ (.A(_19672_),
    .B(_05272_),
    .Y(_05461_));
 sky130_fd_sc_hd__nand3b_4 _27786_ (.A_N(_05461_),
    .B(_05295_),
    .C(_19924_),
    .Y(_05462_));
 sky130_fd_sc_hd__buf_4 _27787_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05463_));
 sky130_fd_sc_hd__buf_4 _27788_ (.A(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__nand2_4 _27789_ (.A(_19685_),
    .B(_05464_),
    .Y(_05465_));
 sky130_vsdinv _27790_ (.A(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__buf_6 _27791_ (.A(_19922_),
    .X(_05467_));
 sky130_fd_sc_hd__nand2_2 _27792_ (.A(_05211_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__nand2_2 _27793_ (.A(_05461_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand3_2 _27794_ (.A(_05462_),
    .B(_05466_),
    .C(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__a22oi_4 _27795_ (.A1(_05280_),
    .A2(_05359_),
    .B1(_05282_),
    .B2(_19920_),
    .Y(_05471_));
 sky130_fd_sc_hd__nor2_4 _27796_ (.A(_05461_),
    .B(_05468_),
    .Y(_05472_));
 sky130_fd_sc_hd__o21ai_2 _27797_ (.A1(_05471_),
    .A2(_05472_),
    .B1(_05465_),
    .Y(_05473_));
 sky130_fd_sc_hd__o211ai_4 _27798_ (.A1(_05362_),
    .A2(_05460_),
    .B1(_05470_),
    .C1(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__a21oi_2 _27799_ (.A1(_05367_),
    .A2(_05364_),
    .B1(_05362_),
    .Y(_05475_));
 sky130_fd_sc_hd__o21ai_2 _27800_ (.A1(_05471_),
    .A2(_05472_),
    .B1(_05466_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand3_2 _27801_ (.A(_05462_),
    .B(_05465_),
    .C(_05469_),
    .Y(_05477_));
 sky130_fd_sc_hd__nand3_4 _27802_ (.A(_05475_),
    .B(_05476_),
    .C(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__nand2_1 _27803_ (.A(_05474_),
    .B(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__buf_4 _27804_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05480_));
 sky130_fd_sc_hd__buf_6 _27805_ (.A(_05480_),
    .X(_05481_));
 sky130_fd_sc_hd__nand2_2 _27806_ (.A(_19682_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__buf_6 _27807_ (.A(_19912_),
    .X(_05483_));
 sky130_fd_sc_hd__buf_6 _27808_ (.A(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__nand3_4 _27809_ (.A(_05482_),
    .B(_19679_),
    .C(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__buf_6 _27810_ (.A(_19912_),
    .X(_05486_));
 sky130_fd_sc_hd__nand2_2 _27811_ (.A(_05125_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__buf_6 _27812_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05488_));
 sky130_fd_sc_hd__buf_4 _27813_ (.A(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__nand3_4 _27814_ (.A(_05487_),
    .B(_05227_),
    .C(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__clkbuf_8 _27815_ (.A(_05132_),
    .X(_05491_));
 sky130_fd_sc_hd__a21oi_1 _27816_ (.A1(_05485_),
    .A2(_05490_),
    .B1(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hd__buf_8 _27817_ (.A(_05208_),
    .X(_05493_));
 sky130_fd_sc_hd__nand2_1 _27818_ (.A(_19676_),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__and3_1 _27819_ (.A(_05485_),
    .B(_05490_),
    .C(_05494_),
    .X(_05495_));
 sky130_fd_sc_hd__a21o_1 _27820_ (.A1(_05492_),
    .A2(_19918_),
    .B1(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__nand2_1 _27821_ (.A(_05479_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__a21oi_4 _27822_ (.A1(_05485_),
    .A2(_05490_),
    .B1(_05494_),
    .Y(_05498_));
 sky130_fd_sc_hd__nor2_4 _27823_ (.A(_05498_),
    .B(_05495_),
    .Y(_05499_));
 sky130_fd_sc_hd__nand3_2 _27824_ (.A(_05499_),
    .B(_05474_),
    .C(_05478_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand3_4 _27825_ (.A(_05459_),
    .B(_05497_),
    .C(_05500_),
    .Y(_05501_));
 sky130_fd_sc_hd__nand3_2 _27826_ (.A(_05496_),
    .B(_05474_),
    .C(_05478_),
    .Y(_05502_));
 sky130_fd_sc_hd__nand2_1 _27827_ (.A(_05479_),
    .B(_05499_),
    .Y(_05503_));
 sky130_fd_sc_hd__o2111ai_4 _27828_ (.A1(_05458_),
    .A2(_05387_),
    .B1(_05372_),
    .C1(_05502_),
    .D1(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__nor2_4 _27829_ (.A(_05376_),
    .B(_05384_),
    .Y(_05505_));
 sky130_fd_sc_hd__o2bb2ai_4 _27830_ (.A1_N(_05501_),
    .A2_N(_05504_),
    .B1(_05381_),
    .B2(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__nor2_2 _27831_ (.A(_05381_),
    .B(_05505_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand3_4 _27832_ (.A(_05504_),
    .B(_05501_),
    .C(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__nand2_2 _27833_ (.A(_05506_),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__nor2_1 _27834_ (.A(_05457_),
    .B(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__and3_1 _27835_ (.A(_05400_),
    .B(_05402_),
    .C(_05413_),
    .X(_05511_));
 sky130_fd_sc_hd__nand2_2 _27836_ (.A(_05509_),
    .B(_05457_),
    .Y(_05512_));
 sky130_fd_sc_hd__nand2_1 _27837_ (.A(_05511_),
    .B(_05512_),
    .Y(_05513_));
 sky130_vsdinv _27838_ (.A(_05457_),
    .Y(_05514_));
 sky130_fd_sc_hd__nand3_4 _27839_ (.A(_05506_),
    .B(_05508_),
    .C(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__a21o_1 _27840_ (.A1(_05512_),
    .A2(_05515_),
    .B1(_05511_),
    .X(_05516_));
 sky130_fd_sc_hd__o21a_1 _27841_ (.A1(_05510_),
    .A2(_05513_),
    .B1(_05516_),
    .X(_05517_));
 sky130_vsdinv _27842_ (.A(_05393_),
    .Y(_05518_));
 sky130_fd_sc_hd__and2_1 _27843_ (.A(_05398_),
    .B(_05401_),
    .X(_05519_));
 sky130_fd_sc_hd__o21bai_2 _27844_ (.A1(_05518_),
    .A2(_05519_),
    .B1_N(_05423_),
    .Y(_05520_));
 sky130_fd_sc_hd__nor2_1 _27845_ (.A(_05518_),
    .B(_05519_),
    .Y(_05521_));
 sky130_fd_sc_hd__nand2_2 _27846_ (.A(_05424_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__nand3_1 _27847_ (.A(_05517_),
    .B(_05520_),
    .C(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__nand2_1 _27848_ (.A(_05520_),
    .B(_05522_),
    .Y(_05524_));
 sky130_fd_sc_hd__nand3_4 _27849_ (.A(_05511_),
    .B(_05512_),
    .C(_05515_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand2_1 _27850_ (.A(_05516_),
    .B(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_1 _27851_ (.A(_05524_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__nand3b_1 _27852_ (.A_N(_05438_),
    .B(_05523_),
    .C(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_1 _27853_ (.A(_05524_),
    .B(_05517_),
    .Y(_05529_));
 sky130_fd_sc_hd__nand3_2 _27854_ (.A(_05526_),
    .B(_05520_),
    .C(_05522_),
    .Y(_05530_));
 sky130_fd_sc_hd__nand3_1 _27855_ (.A(_05529_),
    .B(_05530_),
    .C(_05438_),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_2 _27856_ (.A(_05528_),
    .B(_05531_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _27857_ (.A(_05432_),
    .B(_05433_),
    .Y(_05533_));
 sky130_fd_sc_hd__nand3b_2 _27858_ (.A_N(_05533_),
    .B(_05345_),
    .C(_05354_),
    .Y(_05534_));
 sky130_fd_sc_hd__nand2_2 _27859_ (.A(_05437_),
    .B(_05534_),
    .Y(_05535_));
 sky130_fd_sc_hd__xor2_1 _27860_ (.A(_05532_),
    .B(_05535_),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_2 _27861_ (.A(_05529_),
    .B(_05530_),
    .Y(_05536_));
 sky130_fd_sc_hd__nor2_2 _27862_ (.A(_05345_),
    .B(_05533_),
    .Y(_05537_));
 sky130_fd_sc_hd__a22oi_4 _27863_ (.A1(_05536_),
    .A2(_05537_),
    .B1(_05535_),
    .B2(_05532_),
    .Y(_05538_));
 sky130_fd_sc_hd__a21o_2 _27864_ (.A1(_05501_),
    .A2(_05508_),
    .B1(_05525_),
    .X(_05539_));
 sky130_fd_sc_hd__nand3_2 _27865_ (.A(_05525_),
    .B(_05501_),
    .C(_05508_),
    .Y(_05540_));
 sky130_fd_sc_hd__nand2_1 _27866_ (.A(_05499_),
    .B(_05478_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand2_1 _27867_ (.A(_05541_),
    .B(_05474_),
    .Y(_05542_));
 sky130_fd_sc_hd__nand2_2 _27868_ (.A(_05118_),
    .B(_05464_),
    .Y(_05543_));
 sky130_fd_sc_hd__nand3_4 _27869_ (.A(_05543_),
    .B(_05161_),
    .C(_05489_),
    .Y(_05544_));
 sky130_fd_sc_hd__buf_6 _27870_ (.A(_05480_),
    .X(_05545_));
 sky130_fd_sc_hd__nand2_2 _27871_ (.A(_05125_),
    .B(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__nand3_4 _27872_ (.A(_05546_),
    .B(_05382_),
    .C(_19907_),
    .Y(_05547_));
 sky130_fd_sc_hd__buf_4 _27873_ (.A(_19913_),
    .X(_05548_));
 sky130_fd_sc_hd__nand2_1 _27874_ (.A(_19676_),
    .B(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__a21oi_4 _27875_ (.A1(_05544_),
    .A2(_05547_),
    .B1(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__buf_4 _27876_ (.A(_05278_),
    .X(_05551_));
 sky130_fd_sc_hd__o211a_2 _27877_ (.A1(_05132_),
    .A2(_05551_),
    .B1(_05544_),
    .C1(_05547_),
    .X(_05552_));
 sky130_fd_sc_hd__buf_6 _27878_ (.A(_05267_),
    .X(_05553_));
 sky130_fd_sc_hd__a22oi_4 _27879_ (.A1(_05284_),
    .A2(_05224_),
    .B1(_05366_),
    .B2(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2_2 _27880_ (.A(_19669_),
    .B(_19919_),
    .Y(_05555_));
 sky130_fd_sc_hd__nand2_2 _27881_ (.A(_05201_),
    .B(_05271_),
    .Y(_05556_));
 sky130_fd_sc_hd__nor2_2 _27882_ (.A(_05555_),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__buf_6 _27883_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05558_));
 sky130_fd_sc_hd__nand2_4 _27884_ (.A(_19685_),
    .B(_05558_),
    .Y(_05559_));
 sky130_vsdinv _27885_ (.A(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__o21ai_2 _27886_ (.A1(_05554_),
    .A2(_05557_),
    .B1(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__buf_8 _27887_ (.A(_05168_),
    .X(_05562_));
 sky130_fd_sc_hd__nand3b_4 _27888_ (.A_N(_05555_),
    .B(_05562_),
    .C(_19917_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2_2 _27889_ (.A(_05555_),
    .B(_05556_),
    .Y(_05564_));
 sky130_fd_sc_hd__nand3_2 _27890_ (.A(_05563_),
    .B(_05559_),
    .C(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__a21oi_2 _27891_ (.A1(_05466_),
    .A2(_05469_),
    .B1(_05472_),
    .Y(_05566_));
 sky130_fd_sc_hd__nand3_4 _27892_ (.A(_05561_),
    .B(_05565_),
    .C(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__o21ai_2 _27893_ (.A1(_05554_),
    .A2(_05557_),
    .B1(_05559_),
    .Y(_05568_));
 sky130_fd_sc_hd__nand3_4 _27894_ (.A(_05563_),
    .B(_05560_),
    .C(_05564_),
    .Y(_05569_));
 sky130_fd_sc_hd__o21ai_2 _27895_ (.A1(_05465_),
    .A2(_05471_),
    .B1(_05462_),
    .Y(_05570_));
 sky130_fd_sc_hd__nand3_4 _27896_ (.A(_05568_),
    .B(_05569_),
    .C(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__nand2_1 _27897_ (.A(_05567_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__o21ai_2 _27898_ (.A1(_05550_),
    .A2(_05552_),
    .B1(_05572_),
    .Y(_05573_));
 sky130_fd_sc_hd__nor2_4 _27899_ (.A(_05550_),
    .B(_05552_),
    .Y(_05574_));
 sky130_fd_sc_hd__nand3_2 _27900_ (.A(_05574_),
    .B(_05567_),
    .C(_05571_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand3_4 _27901_ (.A(_05542_),
    .B(_05573_),
    .C(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__a21boi_2 _27902_ (.A1(_05499_),
    .A2(_05478_),
    .B1_N(_05474_),
    .Y(_05577_));
 sky130_fd_sc_hd__nand2_1 _27903_ (.A(_05572_),
    .B(_05574_),
    .Y(_05578_));
 sky130_fd_sc_hd__nand3b_2 _27904_ (.A_N(_05574_),
    .B(_05571_),
    .C(_05567_),
    .Y(_05579_));
 sky130_fd_sc_hd__nand3_4 _27905_ (.A(_05577_),
    .B(_05578_),
    .C(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__nor2_1 _27906_ (.A(_05487_),
    .B(_05482_),
    .Y(_05581_));
 sky130_fd_sc_hd__or2_4 _27907_ (.A(_05581_),
    .B(_05498_),
    .X(_05582_));
 sky130_fd_sc_hd__a21o_1 _27908_ (.A1(_05576_),
    .A2(_05580_),
    .B1(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__nand3_2 _27909_ (.A(_05576_),
    .B(_05580_),
    .C(_05582_),
    .Y(_05584_));
 sky130_fd_sc_hd__a21oi_4 _27910_ (.A1(_05448_),
    .A2(_05445_),
    .B1(_05442_),
    .Y(_05585_));
 sky130_fd_sc_hd__buf_6 _27911_ (.A(_05439_),
    .X(_05586_));
 sky130_fd_sc_hd__buf_6 _27912_ (.A(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__buf_6 _27913_ (.A(\pcpi_mul.rs2[7] ),
    .X(_05588_));
 sky130_fd_sc_hd__buf_6 _27914_ (.A(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__a22oi_4 _27915_ (.A1(_05587_),
    .A2(_05123_),
    .B1(_05589_),
    .B2(_05121_),
    .Y(_05590_));
 sky130_fd_sc_hd__clkbuf_8 _27916_ (.A(_05439_),
    .X(_05591_));
 sky130_fd_sc_hd__nand2_2 _27917_ (.A(_05591_),
    .B(_05441_),
    .Y(_05592_));
 sky130_fd_sc_hd__nand2_2 _27918_ (.A(_19664_),
    .B(_05120_),
    .Y(_05593_));
 sky130_fd_sc_hd__nor2_2 _27919_ (.A(_05592_),
    .B(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_2 _27920_ (.A(_05443_),
    .B(_05146_),
    .Y(_05595_));
 sky130_fd_sc_hd__o21ai_2 _27921_ (.A1(_05590_),
    .A2(_05594_),
    .B1(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__or2_1 _27922_ (.A(_05592_),
    .B(_05593_),
    .X(_05597_));
 sky130_vsdinv _27923_ (.A(_05595_),
    .Y(_05598_));
 sky130_fd_sc_hd__nand2_2 _27924_ (.A(_05592_),
    .B(_05593_),
    .Y(_05599_));
 sky130_fd_sc_hd__nand3_2 _27925_ (.A(_05597_),
    .B(_05598_),
    .C(_05599_),
    .Y(_05600_));
 sky130_fd_sc_hd__nand3b_2 _27926_ (.A_N(_05585_),
    .B(_05596_),
    .C(_05600_),
    .Y(_05601_));
 sky130_fd_sc_hd__clkbuf_4 _27927_ (.A(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__nand3_2 _27928_ (.A(_05597_),
    .B(_05595_),
    .C(_05599_),
    .Y(_05603_));
 sky130_fd_sc_hd__o21ai_2 _27929_ (.A1(_05590_),
    .A2(_05594_),
    .B1(_05598_),
    .Y(_05604_));
 sky130_fd_sc_hd__nand3_4 _27930_ (.A(_05603_),
    .B(_05585_),
    .C(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_4 _27931_ (.A(_05602_),
    .B(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__xor2_4 _27932_ (.A(_05456_),
    .B(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__nand3_4 _27933_ (.A(_05583_),
    .B(_05584_),
    .C(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__a21bo_1 _27934_ (.A1(_05576_),
    .A2(_05580_),
    .B1_N(_05582_),
    .X(_05609_));
 sky130_fd_sc_hd__nand3b_4 _27935_ (.A_N(_05582_),
    .B(_05576_),
    .C(_05580_),
    .Y(_05610_));
 sky130_fd_sc_hd__nand3b_4 _27936_ (.A_N(_05607_),
    .B(_05609_),
    .C(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hd__o2bb2ai_2 _27937_ (.A1_N(_05608_),
    .A2_N(_05611_),
    .B1(_05457_),
    .B2(_05509_),
    .Y(_05612_));
 sky130_fd_sc_hd__nand3b_4 _27938_ (.A_N(_05515_),
    .B(_05608_),
    .C(_05611_),
    .Y(_05613_));
 sky130_fd_sc_hd__nand2_2 _27939_ (.A(_05612_),
    .B(_05613_),
    .Y(_05614_));
 sky130_vsdinv _27940_ (.A(_19658_),
    .Y(_05615_));
 sky130_fd_sc_hd__clkbuf_4 _27941_ (.A(_05615_),
    .X(_05616_));
 sky130_fd_sc_hd__nor2_4 _27942_ (.A(net450),
    .B(_04842_),
    .Y(_05617_));
 sky130_vsdinv _27943_ (.A(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_2 _27944_ (.A(_05614_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__nand3_4 _27945_ (.A(_05612_),
    .B(_05613_),
    .C(_05617_),
    .Y(_05620_));
 sky130_fd_sc_hd__a22oi_2 _27946_ (.A1(_05539_),
    .A2(_05540_),
    .B1(_05619_),
    .B2(_05620_),
    .Y(_05621_));
 sky130_vsdinv _27947_ (.A(_05508_),
    .Y(_05622_));
 sky130_fd_sc_hd__nand2_2 _27948_ (.A(_05525_),
    .B(_05501_),
    .Y(_05623_));
 sky130_fd_sc_hd__o2111a_1 _27949_ (.A1(_05622_),
    .A2(_05623_),
    .B1(_05620_),
    .C1(_05539_),
    .D1(_05619_),
    .X(_05624_));
 sky130_fd_sc_hd__nor2_1 _27950_ (.A(_05521_),
    .B(_05424_),
    .Y(_05625_));
 sky130_fd_sc_hd__a31o_1 _27951_ (.A1(_05516_),
    .A2(_05522_),
    .A3(_05525_),
    .B1(_05625_),
    .X(_05626_));
 sky130_vsdinv _27952_ (.A(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__o21ai_2 _27953_ (.A1(_05621_),
    .A2(_05624_),
    .B1(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__a22o_1 _27954_ (.A1(_05539_),
    .A2(_05540_),
    .B1(_05619_),
    .B2(_05620_),
    .X(_05629_));
 sky130_fd_sc_hd__o2111ai_4 _27955_ (.A1(_05622_),
    .A2(_05623_),
    .B1(_05620_),
    .C1(_05539_),
    .D1(_05619_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand3_4 _27956_ (.A(_05629_),
    .B(_05630_),
    .C(_05626_),
    .Y(_05631_));
 sky130_fd_sc_hd__nand2_2 _27957_ (.A(_05536_),
    .B(_05429_),
    .Y(_05632_));
 sky130_fd_sc_hd__a21boi_4 _27958_ (.A1(_05628_),
    .A2(_05631_),
    .B1_N(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__a31o_1 _27959_ (.A1(_05429_),
    .A2(_05536_),
    .A3(_05628_),
    .B1(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__xor2_1 _27960_ (.A(_05538_),
    .B(_05634_),
    .X(_02686_));
 sky130_vsdinv _27961_ (.A(_05628_),
    .Y(_05635_));
 sky130_fd_sc_hd__o22ai_4 _27962_ (.A1(_05632_),
    .A2(_05635_),
    .B1(_05633_),
    .B2(_05538_),
    .Y(_05636_));
 sky130_fd_sc_hd__buf_6 _27963_ (.A(_05277_),
    .X(_05637_));
 sky130_fd_sc_hd__a22oi_4 _27964_ (.A1(_05280_),
    .A2(_05553_),
    .B1(_05358_),
    .B2(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__nand2_2 _27965_ (.A(_05294_),
    .B(_05377_),
    .Y(_05639_));
 sky130_fd_sc_hd__nand2_2 _27966_ (.A(_19672_),
    .B(_05483_),
    .Y(_05640_));
 sky130_fd_sc_hd__nor2_4 _27967_ (.A(_05639_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__buf_2 _27968_ (.A(\pcpi_mul.rs1[10] ),
    .X(_05642_));
 sky130_fd_sc_hd__buf_4 _27969_ (.A(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__nand2_2 _27970_ (.A(_19685_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__clkbuf_2 _27971_ (.A(_05644_),
    .X(_05645_));
 sky130_fd_sc_hd__o21bai_2 _27972_ (.A1(_05638_),
    .A2(_05641_),
    .B1_N(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__buf_4 _27973_ (.A(_05201_),
    .X(_05647_));
 sky130_fd_sc_hd__nand3b_4 _27974_ (.A_N(_05639_),
    .B(_05647_),
    .C(_05548_),
    .Y(_05648_));
 sky130_fd_sc_hd__nand2_2 _27975_ (.A(_05639_),
    .B(_05640_),
    .Y(_05649_));
 sky130_fd_sc_hd__nand3_2 _27976_ (.A(_05648_),
    .B(_05645_),
    .C(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__o21ai_1 _27977_ (.A1(_05555_),
    .A2(_05556_),
    .B1(_05559_),
    .Y(_05651_));
 sky130_fd_sc_hd__nand2_1 _27978_ (.A(_05651_),
    .B(_05564_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand3_4 _27979_ (.A(_05646_),
    .B(_05650_),
    .C(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__o21ai_2 _27980_ (.A1(_05638_),
    .A2(_05641_),
    .B1(_05645_),
    .Y(_05654_));
 sky130_fd_sc_hd__o21ai_4 _27981_ (.A1(_05559_),
    .A2(_05554_),
    .B1(_05563_),
    .Y(_05655_));
 sky130_fd_sc_hd__buf_6 _27982_ (.A(_05379_),
    .X(_05656_));
 sky130_fd_sc_hd__a41oi_2 _27983_ (.A1(_05295_),
    .A2(_05562_),
    .A3(_05656_),
    .A4(_05383_),
    .B1(_05644_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand2_2 _27984_ (.A(_05657_),
    .B(_05649_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand3_4 _27985_ (.A(_05654_),
    .B(_05655_),
    .C(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__buf_4 _27986_ (.A(\pcpi_mul.rs1[8] ),
    .X(_05660_));
 sky130_fd_sc_hd__buf_6 _27987_ (.A(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__a22oi_4 _27988_ (.A1(_05266_),
    .A2(_05661_),
    .B1(_05382_),
    .B2(_19904_),
    .Y(_05662_));
 sky130_fd_sc_hd__inv_8 _27989_ (.A(_05463_),
    .Y(_05663_));
 sky130_fd_sc_hd__nand3_4 _27990_ (.A(_05116_),
    .B(_19681_),
    .C(_05558_),
    .Y(_05664_));
 sky130_fd_sc_hd__nor2_8 _27991_ (.A(_05663_),
    .B(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__buf_6 _27992_ (.A(_05545_),
    .X(_05666_));
 sky130_fd_sc_hd__nand2_2 _27993_ (.A(_19676_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__o21ai_2 _27994_ (.A1(_05662_),
    .A2(_05665_),
    .B1(_05667_),
    .Y(_05668_));
 sky130_fd_sc_hd__buf_1 _27995_ (.A(_05663_),
    .X(_05669_));
 sky130_fd_sc_hd__buf_6 _27996_ (.A(_05131_),
    .X(_05670_));
 sky130_fd_sc_hd__buf_6 _27997_ (.A(_05481_),
    .X(_05671_));
 sky130_fd_sc_hd__buf_6 _27998_ (.A(_05463_),
    .X(_05672_));
 sky130_fd_sc_hd__buf_6 _27999_ (.A(_19903_),
    .X(_05673_));
 sky130_fd_sc_hd__a22o_1 _28000_ (.A1(_05125_),
    .A2(_05672_),
    .B1(_05152_),
    .B2(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__o2111ai_4 _28001_ (.A1(_05669_),
    .A2(_05664_),
    .B1(_05670_),
    .C1(_05671_),
    .D1(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__nand2_4 _28002_ (.A(_05668_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__a21o_1 _28003_ (.A1(_05653_),
    .A2(_05659_),
    .B1(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__a21boi_2 _28004_ (.A1(_05574_),
    .A2(_05567_),
    .B1_N(_05571_),
    .Y(_05678_));
 sky130_fd_sc_hd__nand3_2 _28005_ (.A(_05653_),
    .B(_05659_),
    .C(_05676_),
    .Y(_05679_));
 sky130_fd_sc_hd__nand3_4 _28006_ (.A(_05677_),
    .B(_05678_),
    .C(_05679_),
    .Y(_05680_));
 sky130_vsdinv _28007_ (.A(_05568_),
    .Y(_05681_));
 sky130_fd_sc_hd__nand2_1 _28008_ (.A(_05569_),
    .B(_05570_),
    .Y(_05682_));
 sky130_fd_sc_hd__o2bb2ai_2 _28009_ (.A1_N(_05567_),
    .A2_N(_05574_),
    .B1(_05681_),
    .B2(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hd__nor3_4 _28010_ (.A(_05667_),
    .B(_05662_),
    .C(_05665_),
    .Y(_05684_));
 sky130_fd_sc_hd__o21a_1 _28011_ (.A1(_05662_),
    .A2(_05665_),
    .B1(_05667_),
    .X(_05685_));
 sky130_fd_sc_hd__o2bb2ai_2 _28012_ (.A1_N(_05653_),
    .A2_N(_05659_),
    .B1(_05684_),
    .B2(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__nand3b_2 _28013_ (.A_N(_05676_),
    .B(_05653_),
    .C(_05659_),
    .Y(_05687_));
 sky130_fd_sc_hd__nand3_4 _28014_ (.A(_05683_),
    .B(_05686_),
    .C(_05687_),
    .Y(_05688_));
 sky130_fd_sc_hd__nor2_4 _28015_ (.A(_05546_),
    .B(_05543_),
    .Y(_05689_));
 sky130_fd_sc_hd__nor2_2 _28016_ (.A(_05689_),
    .B(_05550_),
    .Y(_05690_));
 sky130_vsdinv _28017_ (.A(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__a21oi_4 _28018_ (.A1(_05680_),
    .A2(_05688_),
    .B1(_05691_),
    .Y(_05692_));
 sky130_fd_sc_hd__nand3_4 _28019_ (.A(_05680_),
    .B(_05688_),
    .C(_05691_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand2_2 _28020_ (.A(_05586_),
    .B(_05120_),
    .Y(_05694_));
 sky130_fd_sc_hd__buf_4 _28021_ (.A(_19922_),
    .X(_05695_));
 sky130_fd_sc_hd__nand2_2 _28022_ (.A(_05588_),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__nor2_4 _28023_ (.A(_05694_),
    .B(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__and2_1 _28024_ (.A(_05694_),
    .B(_05696_),
    .X(_05698_));
 sky130_fd_sc_hd__buf_6 _28025_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05699_));
 sky130_fd_sc_hd__nand2_2 _28026_ (.A(_05699_),
    .B(_05174_),
    .Y(_05700_));
 sky130_fd_sc_hd__o21ai_4 _28027_ (.A1(_05697_),
    .A2(_05698_),
    .B1(_05700_),
    .Y(_05701_));
 sky130_vsdinv _28028_ (.A(_05700_),
    .Y(_05702_));
 sky130_fd_sc_hd__nand2_2 _28029_ (.A(_05694_),
    .B(_05696_),
    .Y(_05703_));
 sky130_fd_sc_hd__nand3b_4 _28030_ (.A_N(_05697_),
    .B(_05702_),
    .C(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__nand2_1 _28031_ (.A(_05701_),
    .B(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__a21o_2 _28032_ (.A1(_05598_),
    .A2(_05599_),
    .B1(_05594_),
    .X(_05706_));
 sky130_vsdinv _28033_ (.A(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand2_4 _28034_ (.A(_05705_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__nand3_4 _28035_ (.A(_05701_),
    .B(_05704_),
    .C(_05706_),
    .Y(_05709_));
 sky130_fd_sc_hd__nand2_2 _28036_ (.A(_05708_),
    .B(_05709_),
    .Y(_05710_));
 sky130_fd_sc_hd__nand2_1 _28037_ (.A(_05601_),
    .B(_05456_),
    .Y(_05711_));
 sky130_fd_sc_hd__nand3_1 _28038_ (.A(_05710_),
    .B(_05605_),
    .C(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_1 _28039_ (.A(_05600_),
    .B(_05596_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _28040_ (.A(_05454_),
    .B(_05409_),
    .Y(_05714_));
 sky130_fd_sc_hd__nand3b_4 _28041_ (.A_N(_05714_),
    .B(_05449_),
    .C(_05605_),
    .Y(_05715_));
 sky130_fd_sc_hd__o2111ai_4 _28042_ (.A1(_05585_),
    .A2(_05713_),
    .B1(_05708_),
    .C1(_05709_),
    .D1(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__nand2_2 _28043_ (.A(_05712_),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__nand2_2 _28044_ (.A(_05693_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__o2bb2ai_2 _28045_ (.A1_N(_05680_),
    .A2_N(_05688_),
    .B1(_05689_),
    .B2(_05550_),
    .Y(_05719_));
 sky130_fd_sc_hd__clkbuf_4 _28046_ (.A(_05709_),
    .X(_05720_));
 sky130_fd_sc_hd__a22oi_2 _28047_ (.A1(_05708_),
    .A2(_05720_),
    .B1(_05715_),
    .B2(_05602_),
    .Y(_05721_));
 sky130_fd_sc_hd__a21oi_1 _28048_ (.A1(_05711_),
    .A2(_05605_),
    .B1(_05710_),
    .Y(_05722_));
 sky130_fd_sc_hd__nor2_2 _28049_ (.A(_05721_),
    .B(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__nand3_2 _28050_ (.A(_05680_),
    .B(_05688_),
    .C(_05690_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand3_4 _28051_ (.A(_05719_),
    .B(_05723_),
    .C(_05724_),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_2 _28052_ (.A1(_05692_),
    .A2(_05718_),
    .B1(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_2 _28053_ (.A(_05726_),
    .B(_05608_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand2_1 _28054_ (.A(_05609_),
    .B(_05610_),
    .Y(_05728_));
 sky130_fd_sc_hd__o2111ai_4 _28055_ (.A1(_05692_),
    .A2(_05718_),
    .B1(_05607_),
    .C1(_05725_),
    .D1(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__clkbuf_4 _28056_ (.A(_05729_),
    .X(_05730_));
 sky130_fd_sc_hd__buf_4 _28057_ (.A(\pcpi_mul.rs2[9] ),
    .X(_05731_));
 sky130_fd_sc_hd__buf_6 _28058_ (.A(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__nand2_4 _28059_ (.A(_05732_),
    .B(_19931_),
    .Y(_05733_));
 sky130_fd_sc_hd__and3_4 _28060_ (.A(_05733_),
    .B(net457),
    .C(_19934_),
    .X(_05734_));
 sky130_fd_sc_hd__buf_4 _28061_ (.A(\pcpi_mul.rs2[10] ),
    .X(_05735_));
 sky130_fd_sc_hd__buf_8 _28062_ (.A(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__buf_4 _28063_ (.A(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__nand2_2 _28064_ (.A(net448),
    .B(_05406_),
    .Y(_05738_));
 sky130_fd_sc_hd__and3_2 _28065_ (.A(_05738_),
    .B(net456),
    .C(_19931_),
    .X(_05739_));
 sky130_fd_sc_hd__nor2_4 _28066_ (.A(_05734_),
    .B(_05739_),
    .Y(_05740_));
 sky130_vsdinv _28067_ (.A(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__a21oi_4 _28068_ (.A1(_05727_),
    .A2(_05730_),
    .B1(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__nor2_2 _28069_ (.A(_05620_),
    .B(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand3_2 _28070_ (.A(_05727_),
    .B(_05730_),
    .C(_05741_),
    .Y(_05744_));
 sky130_fd_sc_hd__nand2_2 _28071_ (.A(_05743_),
    .B(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__o211a_2 _28072_ (.A1(_05734_),
    .A2(_05739_),
    .B1(_05730_),
    .C1(_05727_),
    .X(_05746_));
 sky130_fd_sc_hd__o22ai_4 _28073_ (.A1(_05618_),
    .A2(_05614_),
    .B1(_05742_),
    .B2(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__a21boi_4 _28074_ (.A1(_05582_),
    .A2(_05580_),
    .B1_N(_05576_),
    .Y(_05748_));
 sky130_fd_sc_hd__nor2_4 _28075_ (.A(_05748_),
    .B(_05613_),
    .Y(_05749_));
 sky130_fd_sc_hd__and2_1 _28076_ (.A(_05613_),
    .B(_05748_),
    .X(_05750_));
 sky130_fd_sc_hd__nor2_4 _28077_ (.A(_05749_),
    .B(_05750_),
    .Y(_05751_));
 sky130_vsdinv _28078_ (.A(_05751_),
    .Y(_05752_));
 sky130_fd_sc_hd__a21o_1 _28079_ (.A1(_05745_),
    .A2(_05747_),
    .B1(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__and2_1 _28080_ (.A(_05630_),
    .B(_05539_),
    .X(_05754_));
 sky130_fd_sc_hd__nand3_2 _28081_ (.A(_05752_),
    .B(_05745_),
    .C(_05747_),
    .Y(_05755_));
 sky130_fd_sc_hd__nand3_4 _28082_ (.A(_05753_),
    .B(_05754_),
    .C(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__a21o_1 _28083_ (.A1(_05745_),
    .A2(_05747_),
    .B1(_05751_),
    .X(_05757_));
 sky130_fd_sc_hd__nand3_2 _28084_ (.A(_05745_),
    .B(_05751_),
    .C(_05747_),
    .Y(_05758_));
 sky130_fd_sc_hd__nand2_1 _28085_ (.A(_05630_),
    .B(_05539_),
    .Y(_05759_));
 sky130_fd_sc_hd__nand3_2 _28086_ (.A(_05757_),
    .B(_05758_),
    .C(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__nand2_1 _28087_ (.A(_05756_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__nand2_2 _28088_ (.A(_05761_),
    .B(_05631_),
    .Y(_05762_));
 sky130_vsdinv _28089_ (.A(_05631_),
    .Y(_05763_));
 sky130_vsdinv _28090_ (.A(_05762_),
    .Y(_05764_));
 sky130_fd_sc_hd__a21oi_1 _28091_ (.A1(_05763_),
    .A2(_05756_),
    .B1(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__nor2_1 _28092_ (.A(_05636_),
    .B(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__a21oi_2 _28093_ (.A1(_05636_),
    .A2(_05762_),
    .B1(_05766_),
    .Y(_02629_));
 sky130_fd_sc_hd__nand2_1 _28094_ (.A(_05757_),
    .B(_05758_),
    .Y(_05767_));
 sky130_fd_sc_hd__buf_6 _28095_ (.A(_05294_),
    .X(_05768_));
 sky130_fd_sc_hd__buf_6 _28096_ (.A(\pcpi_mul.rs1[7] ),
    .X(_05769_));
 sky130_fd_sc_hd__buf_6 _28097_ (.A(_05769_),
    .X(_05770_));
 sky130_fd_sc_hd__a22oi_4 _28098_ (.A1(_05768_),
    .A2(_05484_),
    .B1(_05647_),
    .B2(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__buf_6 _28099_ (.A(_05294_),
    .X(_05772_));
 sky130_fd_sc_hd__and4_4 _28100_ (.A(_05772_),
    .B(_05282_),
    .C(_19910_),
    .D(_05637_),
    .X(_05773_));
 sky130_fd_sc_hd__buf_6 _28101_ (.A(_19897_),
    .X(_05774_));
 sky130_fd_sc_hd__nand2_4 _28102_ (.A(_05171_),
    .B(_05774_),
    .Y(_05775_));
 sky130_vsdinv _28103_ (.A(_05775_),
    .Y(_05776_));
 sky130_fd_sc_hd__o21ai_2 _28104_ (.A1(_05771_),
    .A2(_05773_),
    .B1(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__clkbuf_4 _28105_ (.A(_05294_),
    .X(_05778_));
 sky130_fd_sc_hd__nand2_1 _28106_ (.A(_05778_),
    .B(_05484_),
    .Y(_05779_));
 sky130_fd_sc_hd__buf_8 _28107_ (.A(_05282_),
    .X(_05780_));
 sky130_fd_sc_hd__nand3b_4 _28108_ (.A_N(_05779_),
    .B(_05780_),
    .C(_19911_),
    .Y(_05781_));
 sky130_fd_sc_hd__a22o_2 _28109_ (.A1(_05768_),
    .A2(_05484_),
    .B1(_05647_),
    .B2(_05770_),
    .X(_05782_));
 sky130_fd_sc_hd__nand3_2 _28110_ (.A(_05781_),
    .B(_05775_),
    .C(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__o21ai_1 _28111_ (.A1(_05639_),
    .A2(_05640_),
    .B1(_05645_),
    .Y(_05784_));
 sky130_fd_sc_hd__nand2_1 _28112_ (.A(_05784_),
    .B(_05649_),
    .Y(_05785_));
 sky130_fd_sc_hd__nand3_4 _28113_ (.A(_05777_),
    .B(_05783_),
    .C(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__clkinv_8 _28114_ (.A(_19897_),
    .Y(_05787_));
 sky130_fd_sc_hd__buf_6 _28115_ (.A(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__o22ai_4 _28116_ (.A1(net474),
    .A2(_05788_),
    .B1(_05771_),
    .B2(_05773_),
    .Y(_05789_));
 sky130_fd_sc_hd__o21ai_2 _28117_ (.A1(_05645_),
    .A2(_05638_),
    .B1(_05648_),
    .Y(_05790_));
 sky130_fd_sc_hd__buf_6 _28118_ (.A(_05203_),
    .X(_05791_));
 sky130_fd_sc_hd__buf_6 _28119_ (.A(_05366_),
    .X(_05792_));
 sky130_fd_sc_hd__a41oi_4 _28120_ (.A1(_05791_),
    .A2(_05792_),
    .A3(_05671_),
    .A4(_19914_),
    .B1(_05775_),
    .Y(_05793_));
 sky130_fd_sc_hd__nand2_2 _28121_ (.A(_05793_),
    .B(_05782_),
    .Y(_05794_));
 sky130_fd_sc_hd__nand3_4 _28122_ (.A(_05789_),
    .B(_05790_),
    .C(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__buf_4 _28123_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05796_));
 sky130_fd_sc_hd__buf_6 _28124_ (.A(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__buf_4 _28125_ (.A(_05642_),
    .X(_05798_));
 sky130_fd_sc_hd__buf_6 _28126_ (.A(_05798_),
    .X(_05799_));
 sky130_fd_sc_hd__a22oi_4 _28127_ (.A1(_05126_),
    .A2(_05797_),
    .B1(_05223_),
    .B2(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__clkbuf_8 _28128_ (.A(\pcpi_mul.rs1[9] ),
    .X(_05801_));
 sky130_fd_sc_hd__clkinv_8 _28129_ (.A(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__buf_2 _28130_ (.A(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__buf_6 _28131_ (.A(_05643_),
    .X(_05804_));
 sky130_fd_sc_hd__nand3_4 _28132_ (.A(_05233_),
    .B(_05382_),
    .C(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__nor2_8 _28133_ (.A(net447),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__buf_6 _28134_ (.A(_19676_),
    .X(_05807_));
 sky130_fd_sc_hd__buf_6 _28135_ (.A(_05661_),
    .X(_05808_));
 sky130_fd_sc_hd__nand2_2 _28136_ (.A(_05807_),
    .B(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__o21ai_1 _28137_ (.A1(_05800_),
    .A2(_05806_),
    .B1(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hd__buf_6 _28138_ (.A(_05643_),
    .X(_05811_));
 sky130_fd_sc_hd__a22o_1 _28139_ (.A1(_05126_),
    .A2(_05797_),
    .B1(_19683_),
    .B2(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__o2111ai_4 _28140_ (.A1(net447),
    .A2(_05805_),
    .B1(_19677_),
    .C1(_19908_),
    .D1(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__nand2_2 _28141_ (.A(_05810_),
    .B(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__a21o_1 _28142_ (.A1(_05786_),
    .A2(_05795_),
    .B1(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__nand2_1 _28143_ (.A(_05659_),
    .B(_05676_),
    .Y(_05816_));
 sky130_fd_sc_hd__nand2_1 _28144_ (.A(_05816_),
    .B(_05653_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand3_2 _28145_ (.A(_05786_),
    .B(_05795_),
    .C(_05814_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand3_4 _28146_ (.A(_05815_),
    .B(_05817_),
    .C(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__o21a_1 _28147_ (.A1(_05638_),
    .A2(_05641_),
    .B1(_05645_),
    .X(_05820_));
 sky130_fd_sc_hd__nand2_1 _28148_ (.A(_05655_),
    .B(_05658_),
    .Y(_05821_));
 sky130_fd_sc_hd__a21oi_2 _28149_ (.A1(_05654_),
    .A2(_05658_),
    .B1(_05655_),
    .Y(_05822_));
 sky130_fd_sc_hd__o22ai_4 _28150_ (.A1(_05820_),
    .A2(_05821_),
    .B1(_05676_),
    .B2(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__nor3_4 _28151_ (.A(_05809_),
    .B(_05800_),
    .C(_05806_),
    .Y(_05824_));
 sky130_fd_sc_hd__o21a_1 _28152_ (.A1(_05800_),
    .A2(_05806_),
    .B1(_05809_),
    .X(_05825_));
 sky130_fd_sc_hd__o2bb2ai_2 _28153_ (.A1_N(_05795_),
    .A2_N(_05786_),
    .B1(_05824_),
    .B2(_05825_),
    .Y(_05826_));
 sky130_fd_sc_hd__nand3b_2 _28154_ (.A_N(_05814_),
    .B(_05786_),
    .C(_05795_),
    .Y(_05827_));
 sky130_fd_sc_hd__nand3_4 _28155_ (.A(_05823_),
    .B(_05826_),
    .C(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__nor2_1 _28156_ (.A(_05665_),
    .B(_05684_),
    .Y(_05829_));
 sky130_vsdinv _28157_ (.A(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__a21o_1 _28158_ (.A1(_05819_),
    .A2(_05828_),
    .B1(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__buf_6 _28159_ (.A(_05450_),
    .X(_05832_));
 sky130_fd_sc_hd__buf_6 _28160_ (.A(_05403_),
    .X(_05833_));
 sky130_fd_sc_hd__nand3_4 _28161_ (.A(_05832_),
    .B(_05833_),
    .C(_05374_),
    .Y(_05834_));
 sky130_fd_sc_hd__buf_6 _28162_ (.A(\pcpi_mul.rs2[6] ),
    .X(_05835_));
 sky130_fd_sc_hd__nand2_2 _28163_ (.A(_05835_),
    .B(_05383_),
    .Y(_05836_));
 sky130_fd_sc_hd__buf_6 _28164_ (.A(_05591_),
    .X(_05837_));
 sky130_fd_sc_hd__buf_6 _28165_ (.A(_05695_),
    .X(_05838_));
 sky130_fd_sc_hd__a22o_2 _28166_ (.A1(_05837_),
    .A2(_05838_),
    .B1(_19665_),
    .B2(_05225_),
    .X(_05839_));
 sky130_fd_sc_hd__o211ai_4 _28167_ (.A1(_05155_),
    .A2(_05834_),
    .B1(_05836_),
    .C1(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__buf_6 _28168_ (.A(_19661_),
    .X(_05841_));
 sky130_fd_sc_hd__buf_4 _28169_ (.A(_05403_),
    .X(_05842_));
 sky130_fd_sc_hd__buf_6 _28170_ (.A(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__a22oi_4 _28171_ (.A1(_05841_),
    .A2(_05147_),
    .B1(_05843_),
    .B2(_05225_),
    .Y(_05844_));
 sky130_fd_sc_hd__nor2_2 _28172_ (.A(_05155_),
    .B(_05834_),
    .Y(_05845_));
 sky130_vsdinv _28173_ (.A(_05836_),
    .Y(_05846_));
 sky130_fd_sc_hd__o21ai_2 _28174_ (.A1(_05844_),
    .A2(_05845_),
    .B1(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hd__o211ai_4 _28175_ (.A1(_05738_),
    .A2(_05733_),
    .B1(_05840_),
    .C1(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__o21ai_2 _28176_ (.A1(_05844_),
    .A2(_05845_),
    .B1(_05836_),
    .Y(_05849_));
 sky130_fd_sc_hd__nor2_2 _28177_ (.A(_05738_),
    .B(_05733_),
    .Y(_05850_));
 sky130_fd_sc_hd__o211ai_2 _28178_ (.A1(_05155_),
    .A2(_05834_),
    .B1(_05846_),
    .C1(_05839_),
    .Y(_05851_));
 sky130_fd_sc_hd__nand3_4 _28179_ (.A(_05849_),
    .B(_05850_),
    .C(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__a31o_2 _28180_ (.A1(_05703_),
    .A2(_19668_),
    .A3(_19921_),
    .B1(_05697_),
    .X(_05853_));
 sky130_fd_sc_hd__a21o_2 _28181_ (.A1(_05848_),
    .A2(_05852_),
    .B1(_05853_),
    .X(_05854_));
 sky130_fd_sc_hd__nand3_4 _28182_ (.A(_05848_),
    .B(_05852_),
    .C(_05853_),
    .Y(_05855_));
 sky130_fd_sc_hd__nand2_4 _28183_ (.A(_05854_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__a21oi_4 _28184_ (.A1(_05701_),
    .A2(_05704_),
    .B1(_05706_),
    .Y(_05857_));
 sky130_fd_sc_hd__o21ai_1 _28185_ (.A1(_05602_),
    .A2(_05857_),
    .B1(_05720_),
    .Y(_05858_));
 sky130_fd_sc_hd__nand2_1 _28186_ (.A(_05856_),
    .B(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__o2111ai_4 _28187_ (.A1(_05602_),
    .A2(_05857_),
    .B1(_05720_),
    .C1(_05855_),
    .D1(_05854_),
    .Y(_05860_));
 sky130_fd_sc_hd__nand2_1 _28188_ (.A(_05859_),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__nand3_2 _28189_ (.A(_05819_),
    .B(_05828_),
    .C(_05830_),
    .Y(_05862_));
 sky130_fd_sc_hd__nand3_4 _28190_ (.A(_05831_),
    .B(_05861_),
    .C(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__o2bb2ai_2 _28191_ (.A1_N(_05819_),
    .A2_N(_05828_),
    .B1(_05665_),
    .B2(_05684_),
    .Y(_05864_));
 sky130_fd_sc_hd__nand2_1 _28192_ (.A(_05602_),
    .B(_05720_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21oi_1 _28193_ (.A1(_05848_),
    .A2(_05852_),
    .B1(_05853_),
    .Y(_05866_));
 sky130_vsdinv _28194_ (.A(_05855_),
    .Y(_05867_));
 sky130_fd_sc_hd__o2bb2ai_1 _28195_ (.A1_N(_05708_),
    .A2_N(_05865_),
    .B1(_05866_),
    .B2(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__nand3_1 _28196_ (.A(_05858_),
    .B(_05855_),
    .C(_05854_),
    .Y(_05869_));
 sky130_fd_sc_hd__nand2_1 _28197_ (.A(_05868_),
    .B(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__nand3_2 _28198_ (.A(_05819_),
    .B(_05828_),
    .C(_05829_),
    .Y(_05871_));
 sky130_fd_sc_hd__nand3_4 _28199_ (.A(_05864_),
    .B(_05870_),
    .C(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand2_1 _28200_ (.A(_05863_),
    .B(_05872_),
    .Y(_05873_));
 sky130_fd_sc_hd__nand2_1 _28201_ (.A(_05680_),
    .B(_05688_),
    .Y(_05874_));
 sky130_fd_sc_hd__nand2_1 _28202_ (.A(_05874_),
    .B(_05690_),
    .Y(_05875_));
 sky130_fd_sc_hd__nor3_4 _28203_ (.A(_05456_),
    .B(_05606_),
    .C(_05710_),
    .Y(_05876_));
 sky130_fd_sc_hd__a31oi_4 _28204_ (.A1(_05875_),
    .A2(_05717_),
    .A3(_05693_),
    .B1(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__nand2_4 _28205_ (.A(_05873_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__o21bai_2 _28206_ (.A1(_05692_),
    .A2(_05718_),
    .B1_N(_05876_),
    .Y(_05879_));
 sky130_fd_sc_hd__nand3_4 _28207_ (.A(_05879_),
    .B(_05872_),
    .C(_05863_),
    .Y(_05880_));
 sky130_fd_sc_hd__nor2_8 _28208_ (.A(net450),
    .B(_05151_),
    .Y(_05881_));
 sky130_fd_sc_hd__buf_6 _28209_ (.A(\pcpi_mul.rs2[10] ),
    .X(_05882_));
 sky130_fd_sc_hd__buf_8 _28210_ (.A(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__nand2_2 _28211_ (.A(_05883_),
    .B(_05123_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand2_1 _28212_ (.A(net477),
    .B(_05213_),
    .Y(_05885_));
 sky130_fd_sc_hd__nor2_2 _28213_ (.A(_05884_),
    .B(_05885_),
    .Y(_05886_));
 sky130_vsdinv _28214_ (.A(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__nand2_2 _28215_ (.A(_05884_),
    .B(_05885_),
    .Y(_05888_));
 sky130_fd_sc_hd__nand2_2 _28216_ (.A(_05887_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__nor2_2 _28217_ (.A(_05881_),
    .B(_05889_),
    .Y(_05890_));
 sky130_fd_sc_hd__and2_1 _28218_ (.A(_05889_),
    .B(_05881_),
    .X(_05891_));
 sky130_fd_sc_hd__nor2_1 _28219_ (.A(_05890_),
    .B(_05891_),
    .Y(_05892_));
 sky130_vsdinv _28220_ (.A(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__a21o_1 _28221_ (.A1(_05878_),
    .A2(_05880_),
    .B1(_05893_),
    .X(_05894_));
 sky130_fd_sc_hd__nand3_2 _28222_ (.A(_05878_),
    .B(_05880_),
    .C(_05893_),
    .Y(_05895_));
 sky130_fd_sc_hd__nand3_4 _28223_ (.A(_05894_),
    .B(_05746_),
    .C(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__nand2_1 _28224_ (.A(_05727_),
    .B(_05730_),
    .Y(_05897_));
 sky130_fd_sc_hd__a21oi_2 _28225_ (.A1(_05878_),
    .A2(_05880_),
    .B1(_05893_),
    .Y(_05898_));
 sky130_fd_sc_hd__o211a_4 _28226_ (.A1(_05891_),
    .A2(_05890_),
    .B1(_05880_),
    .C1(_05878_),
    .X(_05899_));
 sky130_fd_sc_hd__o22ai_4 _28227_ (.A1(_05740_),
    .A2(_05897_),
    .B1(_05898_),
    .B2(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__and2_2 _28228_ (.A(_05693_),
    .B(_05688_),
    .X(_05901_));
 sky130_fd_sc_hd__nor2_1 _28229_ (.A(_05608_),
    .B(_05726_),
    .Y(_05902_));
 sky130_fd_sc_hd__nor2_1 _28230_ (.A(_05901_),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__and2_1 _28231_ (.A(_05902_),
    .B(_05901_),
    .X(_05904_));
 sky130_fd_sc_hd__o2bb2ai_1 _28232_ (.A1_N(_05896_),
    .A2_N(_05900_),
    .B1(_05903_),
    .B2(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__a22oi_2 _28233_ (.A1(_05743_),
    .A2(_05744_),
    .B1(_05747_),
    .B2(_05751_),
    .Y(_05906_));
 sky130_fd_sc_hd__nor2_4 _28234_ (.A(_05901_),
    .B(_05730_),
    .Y(_05907_));
 sky130_fd_sc_hd__and2_1 _28235_ (.A(_05729_),
    .B(_05901_),
    .X(_05908_));
 sky130_fd_sc_hd__nor2_2 _28236_ (.A(_05907_),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__nand3b_2 _28237_ (.A_N(_05909_),
    .B(_05900_),
    .C(_05896_),
    .Y(_05910_));
 sky130_fd_sc_hd__nand3_2 _28238_ (.A(_05905_),
    .B(_05906_),
    .C(_05910_),
    .Y(_05911_));
 sky130_fd_sc_hd__and2_1 _28239_ (.A(_05911_),
    .B(_05749_),
    .X(_05912_));
 sky130_fd_sc_hd__a21o_1 _28240_ (.A1(_05900_),
    .A2(_05896_),
    .B1(_05909_),
    .X(_05913_));
 sky130_fd_sc_hd__nand2_1 _28241_ (.A(_05747_),
    .B(_05751_),
    .Y(_05914_));
 sky130_fd_sc_hd__nand2_1 _28242_ (.A(_05914_),
    .B(_05745_),
    .Y(_05915_));
 sky130_fd_sc_hd__nand3_1 _28243_ (.A(_05900_),
    .B(_05896_),
    .C(_05909_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand3_2 _28244_ (.A(_05913_),
    .B(_05915_),
    .C(_05916_),
    .Y(_05917_));
 sky130_fd_sc_hd__a21oi_1 _28245_ (.A1(_05917_),
    .A2(_05911_),
    .B1(_05749_),
    .Y(_05918_));
 sky130_fd_sc_hd__o22ai_1 _28246_ (.A1(_05754_),
    .A2(_05767_),
    .B1(_05912_),
    .B2(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__a21o_1 _28247_ (.A1(_05917_),
    .A2(_05911_),
    .B1(_05749_),
    .X(_05920_));
 sky130_vsdinv _28248_ (.A(_05760_),
    .Y(_05921_));
 sky130_fd_sc_hd__nand2_1 _28249_ (.A(_05911_),
    .B(_05749_),
    .Y(_05922_));
 sky130_fd_sc_hd__nand3_1 _28250_ (.A(_05920_),
    .B(_05921_),
    .C(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__nand2_2 _28251_ (.A(_05919_),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__a22oi_4 _28252_ (.A1(_05763_),
    .A2(_05756_),
    .B1(_05636_),
    .B2(_05762_),
    .Y(_05925_));
 sky130_fd_sc_hd__xor2_1 _28253_ (.A(_05924_),
    .B(_05925_),
    .X(_02630_));
 sky130_fd_sc_hd__a21oi_4 _28254_ (.A1(_05881_),
    .A2(_05888_),
    .B1(_05886_),
    .Y(_05926_));
 sky130_fd_sc_hd__nand2_4 _28255_ (.A(_05832_),
    .B(_05374_),
    .Y(_05927_));
 sky130_fd_sc_hd__nand2_4 _28256_ (.A(_05833_),
    .B(_05383_),
    .Y(_05928_));
 sky130_fd_sc_hd__nor2_8 _28257_ (.A(_05927_),
    .B(_05928_),
    .Y(_05929_));
 sky130_vsdinv _28258_ (.A(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__nand2_2 _28259_ (.A(_05699_),
    .B(_05548_),
    .Y(_05931_));
 sky130_vsdinv _28260_ (.A(_05931_),
    .Y(_05932_));
 sky130_fd_sc_hd__nand2_1 _28261_ (.A(_05927_),
    .B(_05928_),
    .Y(_05933_));
 sky130_fd_sc_hd__nand3_2 _28262_ (.A(_05930_),
    .B(_05932_),
    .C(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__and2_2 _28263_ (.A(_05927_),
    .B(_05928_),
    .X(_05935_));
 sky130_fd_sc_hd__o21ai_2 _28264_ (.A1(_05929_),
    .A2(_05935_),
    .B1(_05931_),
    .Y(_05936_));
 sky130_fd_sc_hd__nand3b_4 _28265_ (.A_N(_05926_),
    .B(_05934_),
    .C(_05936_),
    .Y(_05937_));
 sky130_fd_sc_hd__nand3_2 _28266_ (.A(_05930_),
    .B(_05931_),
    .C(_05933_),
    .Y(_05938_));
 sky130_fd_sc_hd__o21ai_2 _28267_ (.A1(_05929_),
    .A2(_05935_),
    .B1(_05932_),
    .Y(_05939_));
 sky130_fd_sc_hd__nand3_4 _28268_ (.A(_05938_),
    .B(_05939_),
    .C(_05926_),
    .Y(_05940_));
 sky130_fd_sc_hd__o21a_2 _28269_ (.A1(_05846_),
    .A2(_05845_),
    .B1(_05839_),
    .X(_05941_));
 sky130_fd_sc_hd__a21o_1 _28270_ (.A1(_05937_),
    .A2(_05940_),
    .B1(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__nand3_4 _28271_ (.A(_05937_),
    .B(_05940_),
    .C(_05941_),
    .Y(_05943_));
 sky130_fd_sc_hd__nand2_2 _28272_ (.A(_05942_),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__nand2_1 _28273_ (.A(_05848_),
    .B(_05853_),
    .Y(_05945_));
 sky130_fd_sc_hd__nand2_2 _28274_ (.A(_05945_),
    .B(_05852_),
    .Y(_05946_));
 sky130_vsdinv _28275_ (.A(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__nand2_1 _28276_ (.A(_05944_),
    .B(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__nor2_2 _28277_ (.A(_05720_),
    .B(_05856_),
    .Y(_05949_));
 sky130_fd_sc_hd__nand3_2 _28278_ (.A(_05942_),
    .B(_05943_),
    .C(_05946_),
    .Y(_05950_));
 sky130_fd_sc_hd__nand3_4 _28279_ (.A(_05948_),
    .B(_05949_),
    .C(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__a21oi_2 _28280_ (.A1(_05942_),
    .A2(_05943_),
    .B1(_05946_),
    .Y(_05952_));
 sky130_fd_sc_hd__and3_4 _28281_ (.A(_05942_),
    .B(_05943_),
    .C(_05946_),
    .X(_05953_));
 sky130_fd_sc_hd__o22ai_4 _28282_ (.A1(_05720_),
    .A2(_05856_),
    .B1(_05952_),
    .B2(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__a21oi_2 _28283_ (.A1(_05789_),
    .A2(_05794_),
    .B1(_05790_),
    .Y(_05955_));
 sky130_fd_sc_hd__o21ai_4 _28284_ (.A1(_05814_),
    .A2(_05955_),
    .B1(_05795_),
    .Y(_05956_));
 sky130_fd_sc_hd__nand2_4 _28285_ (.A(_05295_),
    .B(_19910_),
    .Y(_05957_));
 sky130_fd_sc_hd__buf_6 _28286_ (.A(_05660_),
    .X(_05958_));
 sky130_fd_sc_hd__nand2_4 _28287_ (.A(_05562_),
    .B(_05958_),
    .Y(_05959_));
 sky130_fd_sc_hd__nor2_8 _28288_ (.A(_05957_),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__and2_1 _28289_ (.A(_05957_),
    .B(_05959_),
    .X(_05961_));
 sky130_fd_sc_hd__buf_6 _28290_ (.A(_19893_),
    .X(_05962_));
 sky130_fd_sc_hd__nand2_2 _28291_ (.A(_05171_),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__o21ai_2 _28292_ (.A1(_05960_),
    .A2(_05961_),
    .B1(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__or2_2 _28293_ (.A(_05957_),
    .B(_05959_),
    .X(_05965_));
 sky130_vsdinv _28294_ (.A(_05963_),
    .Y(_05966_));
 sky130_fd_sc_hd__nand2_4 _28295_ (.A(_05957_),
    .B(_05959_),
    .Y(_05967_));
 sky130_fd_sc_hd__nand3_4 _28296_ (.A(_05965_),
    .B(_05966_),
    .C(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__o21ai_4 _28297_ (.A1(_05775_),
    .A2(_05771_),
    .B1(_05781_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand3_4 _28298_ (.A(_05964_),
    .B(_05968_),
    .C(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__o21ai_2 _28299_ (.A1(_05960_),
    .A2(_05961_),
    .B1(_05966_),
    .Y(_05971_));
 sky130_fd_sc_hd__nand3_2 _28300_ (.A(_05965_),
    .B(_05963_),
    .C(_05967_),
    .Y(_05972_));
 sky130_fd_sc_hd__a21oi_4 _28301_ (.A1(_05782_),
    .A2(_05776_),
    .B1(_05773_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand3_4 _28302_ (.A(_05971_),
    .B(_05972_),
    .C(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__nand2_1 _28303_ (.A(_05970_),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__buf_4 _28304_ (.A(\pcpi_mul.rs1[11] ),
    .X(_05976_));
 sky130_fd_sc_hd__buf_6 _28305_ (.A(_05976_),
    .X(_05977_));
 sky130_fd_sc_hd__and4_2 _28306_ (.A(_05117_),
    .B(_05119_),
    .C(_05977_),
    .D(_05811_),
    .X(_05978_));
 sky130_fd_sc_hd__nand2_1 _28307_ (.A(_05162_),
    .B(_19902_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21a_1 _28308_ (.A1(_05153_),
    .A2(_05788_),
    .B1(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__buf_6 _28309_ (.A(_05802_),
    .X(_05981_));
 sky130_fd_sc_hd__nor2_2 _28310_ (.A(_05491_),
    .B(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__o21bai_2 _28311_ (.A1(_05978_),
    .A2(_05980_),
    .B1_N(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__o21ai_2 _28312_ (.A1(_05153_),
    .A2(_05788_),
    .B1(_05979_),
    .Y(_05984_));
 sky130_fd_sc_hd__nand3b_4 _28313_ (.A_N(_05978_),
    .B(_05982_),
    .C(_05984_),
    .Y(_05985_));
 sky130_fd_sc_hd__and2_1 _28314_ (.A(_05983_),
    .B(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__nand2_1 _28315_ (.A(_05975_),
    .B(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__nand2_2 _28316_ (.A(_05983_),
    .B(_05985_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand3_2 _28317_ (.A(_05974_),
    .B(_05988_),
    .C(_05970_),
    .Y(_05989_));
 sky130_fd_sc_hd__nand3b_4 _28318_ (.A_N(_05956_),
    .B(_05987_),
    .C(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__nand2_2 _28319_ (.A(_05975_),
    .B(_05988_),
    .Y(_05991_));
 sky130_fd_sc_hd__nand3_4 _28320_ (.A(_05986_),
    .B(_05974_),
    .C(_05970_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand3_4 _28321_ (.A(_05991_),
    .B(_05992_),
    .C(_05956_),
    .Y(_05993_));
 sky130_fd_sc_hd__nor2_4 _28322_ (.A(_05806_),
    .B(_05824_),
    .Y(_05994_));
 sky130_vsdinv _28323_ (.A(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__a21oi_2 _28324_ (.A1(_05990_),
    .A2(_05993_),
    .B1(_05995_),
    .Y(_05996_));
 sky130_fd_sc_hd__and3_2 _28325_ (.A(_05991_),
    .B(_05992_),
    .C(_05956_),
    .X(_05997_));
 sky130_fd_sc_hd__nand2_2 _28326_ (.A(_05990_),
    .B(_05995_),
    .Y(_05998_));
 sky130_fd_sc_hd__nor2_2 _28327_ (.A(_05997_),
    .B(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__o2bb2ai_2 _28328_ (.A1_N(_05951_),
    .A2_N(_05954_),
    .B1(_05996_),
    .B2(_05999_),
    .Y(_06000_));
 sky130_fd_sc_hd__or2_1 _28329_ (.A(_05602_),
    .B(_05710_),
    .X(_06001_));
 sky130_fd_sc_hd__o21ai_2 _28330_ (.A1(_05856_),
    .A2(_06001_),
    .B1(_05863_),
    .Y(_06002_));
 sky130_fd_sc_hd__nand2_1 _28331_ (.A(_05990_),
    .B(_05993_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand2_1 _28332_ (.A(_06003_),
    .B(_05994_),
    .Y(_06004_));
 sky130_fd_sc_hd__o2111ai_4 _28333_ (.A1(_05997_),
    .A2(_05998_),
    .B1(_05951_),
    .C1(_06004_),
    .D1(_05954_),
    .Y(_06005_));
 sky130_fd_sc_hd__nand3_4 _28334_ (.A(_06000_),
    .B(_06002_),
    .C(_06005_),
    .Y(_06006_));
 sky130_fd_sc_hd__o211ai_2 _28335_ (.A1(_05996_),
    .A2(_05999_),
    .B1(_05954_),
    .C1(_05951_),
    .Y(_06007_));
 sky130_fd_sc_hd__a21oi_1 _28336_ (.A1(_05990_),
    .A2(_05993_),
    .B1(_05994_),
    .Y(_06008_));
 sky130_fd_sc_hd__nor2_1 _28337_ (.A(_05995_),
    .B(_06003_),
    .Y(_06009_));
 sky130_fd_sc_hd__o2bb2ai_2 _28338_ (.A1_N(_05951_),
    .A2_N(_05954_),
    .B1(_06008_),
    .B2(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__o21a_1 _28339_ (.A1(_05856_),
    .A2(_06001_),
    .B1(_05863_),
    .X(_06011_));
 sky130_fd_sc_hd__nand3_4 _28340_ (.A(_06007_),
    .B(_06010_),
    .C(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__buf_6 _28341_ (.A(\pcpi_mul.rs2[9] ),
    .X(_06013_));
 sky130_fd_sc_hd__buf_8 _28342_ (.A(_06013_),
    .X(_06014_));
 sky130_fd_sc_hd__buf_6 _28343_ (.A(_05359_),
    .X(_06015_));
 sky130_fd_sc_hd__nand2_2 _28344_ (.A(_06014_),
    .B(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__buf_2 _28345_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06017_));
 sky130_fd_sc_hd__clkbuf_8 _28346_ (.A(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__buf_8 _28347_ (.A(_05735_),
    .X(_06019_));
 sky130_fd_sc_hd__buf_6 _28348_ (.A(_05229_),
    .X(_06020_));
 sky130_fd_sc_hd__a22oi_4 _28349_ (.A1(_06018_),
    .A2(_05199_),
    .B1(_06019_),
    .B2(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__buf_4 _28350_ (.A(_06017_),
    .X(_06022_));
 sky130_fd_sc_hd__nand2_2 _28351_ (.A(_06022_),
    .B(_19930_),
    .Y(_06023_));
 sky130_fd_sc_hd__buf_6 _28352_ (.A(\pcpi_mul.rs2[10] ),
    .X(_06024_));
 sky130_fd_sc_hd__nand2_2 _28353_ (.A(_06024_),
    .B(_19927_),
    .Y(_06025_));
 sky130_fd_sc_hd__nor2_4 _28354_ (.A(_06023_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__nor3_2 _28355_ (.A(_06016_),
    .B(_06021_),
    .C(_06026_),
    .Y(_06027_));
 sky130_vsdinv _28356_ (.A(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__o21ai_2 _28357_ (.A1(_06021_),
    .A2(_06026_),
    .B1(_06016_),
    .Y(_06029_));
 sky130_vsdinv _28358_ (.A(\pcpi_mul.rs2[12] ),
    .Y(_06030_));
 sky130_fd_sc_hd__clkbuf_4 _28359_ (.A(_06030_),
    .X(_06031_));
 sky130_fd_sc_hd__nor2_8 _28360_ (.A(_06031_),
    .B(net453),
    .Y(_06032_));
 sky130_fd_sc_hd__a21oi_4 _28361_ (.A1(_06028_),
    .A2(_06029_),
    .B1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__and3b_1 _28362_ (.A_N(_06027_),
    .B(_06032_),
    .C(_06029_),
    .X(_06034_));
 sky130_fd_sc_hd__clkbuf_4 _28363_ (.A(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__o2bb2ai_4 _28364_ (.A1_N(_06006_),
    .A2_N(_06012_),
    .B1(_06033_),
    .B2(_06035_),
    .Y(_06036_));
 sky130_fd_sc_hd__nor2_2 _28365_ (.A(_06033_),
    .B(_06035_),
    .Y(_06037_));
 sky130_fd_sc_hd__nand3_4 _28366_ (.A(_06012_),
    .B(_06006_),
    .C(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__a21oi_4 _28367_ (.A1(_06036_),
    .A2(_06038_),
    .B1(_05899_),
    .Y(_06039_));
 sky130_fd_sc_hd__and3_1 _28368_ (.A(_06036_),
    .B(_05899_),
    .C(_06038_),
    .X(_06040_));
 sky130_vsdinv _28369_ (.A(_05828_),
    .Y(_06041_));
 sky130_fd_sc_hd__a21oi_4 _28370_ (.A1(_05830_),
    .A2(_05819_),
    .B1(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__nor2_8 _28371_ (.A(_06042_),
    .B(_05880_),
    .Y(_06043_));
 sky130_fd_sc_hd__and2_1 _28372_ (.A(_05880_),
    .B(_06042_),
    .X(_06044_));
 sky130_fd_sc_hd__nor2_4 _28373_ (.A(_06043_),
    .B(_06044_),
    .Y(_06045_));
 sky130_fd_sc_hd__o21ai_2 _28374_ (.A1(_06039_),
    .A2(_06040_),
    .B1(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__nand2_1 _28375_ (.A(_05900_),
    .B(_05909_),
    .Y(_06047_));
 sky130_fd_sc_hd__and2_1 _28376_ (.A(_06047_),
    .B(_05896_),
    .X(_06048_));
 sky130_fd_sc_hd__a21o_1 _28377_ (.A1(_06036_),
    .A2(_06038_),
    .B1(_05899_),
    .X(_06049_));
 sky130_vsdinv _28378_ (.A(_06045_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand3_2 _28379_ (.A(_06036_),
    .B(_05899_),
    .C(_06038_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand3_2 _28380_ (.A(_06049_),
    .B(_06050_),
    .C(_06051_),
    .Y(_06052_));
 sky130_fd_sc_hd__nand3_4 _28381_ (.A(_06046_),
    .B(_06048_),
    .C(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__nand2_4 _28382_ (.A(_06053_),
    .B(_05907_),
    .Y(_06054_));
 sky130_fd_sc_hd__o22ai_2 _28383_ (.A1(_06043_),
    .A2(_06044_),
    .B1(_06039_),
    .B2(_06040_),
    .Y(_06055_));
 sky130_fd_sc_hd__nand3_1 _28384_ (.A(_06049_),
    .B(_06045_),
    .C(_06051_),
    .Y(_06056_));
 sky130_fd_sc_hd__nand2_1 _28385_ (.A(_06047_),
    .B(_05896_),
    .Y(_06057_));
 sky130_fd_sc_hd__nand3_2 _28386_ (.A(_06055_),
    .B(_06056_),
    .C(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_1 _28387_ (.A(_06053_),
    .B(_06058_),
    .Y(_06059_));
 sky130_vsdinv _28388_ (.A(_05907_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _28389_ (.A(_05922_),
    .B(_05917_),
    .Y(_06061_));
 sky130_fd_sc_hd__a21boi_4 _28390_ (.A1(_06059_),
    .A2(_06060_),
    .B1_N(_06061_),
    .Y(_06062_));
 sky130_fd_sc_hd__o2bb2ai_1 _28391_ (.A1_N(_06058_),
    .A2_N(_06053_),
    .B1(_05730_),
    .B2(_05901_),
    .Y(_06063_));
 sky130_fd_sc_hd__a21oi_2 _28392_ (.A1(_06063_),
    .A2(_06054_),
    .B1(_06061_),
    .Y(_06064_));
 sky130_fd_sc_hd__a21oi_4 _28393_ (.A1(_06054_),
    .A2(_06062_),
    .B1(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_1 _28394_ (.A(_05920_),
    .B(_05921_),
    .Y(_06066_));
 sky130_fd_sc_hd__o22ai_4 _28395_ (.A1(_05912_),
    .A2(_06066_),
    .B1(_05924_),
    .B2(_05925_),
    .Y(_06067_));
 sky130_fd_sc_hd__xor2_1 _28396_ (.A(_06065_),
    .B(_06067_),
    .X(_02631_));
 sky130_fd_sc_hd__nand2_2 _28397_ (.A(_06005_),
    .B(_05951_),
    .Y(_06068_));
 sky130_fd_sc_hd__nor2_2 _28398_ (.A(_06016_),
    .B(_06021_),
    .Y(_06069_));
 sky130_fd_sc_hd__nand3_4 _28399_ (.A(_05832_),
    .B(_05833_),
    .C(_05378_),
    .Y(_06070_));
 sky130_fd_sc_hd__nand2_2 _28400_ (.A(_05835_),
    .B(_19910_),
    .Y(_06071_));
 sky130_vsdinv _28401_ (.A(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__buf_6 _28402_ (.A(_05553_),
    .X(_06073_));
 sky130_fd_sc_hd__a22o_2 _28403_ (.A1(_05841_),
    .A2(_06073_),
    .B1(_05843_),
    .B2(_19914_),
    .X(_06074_));
 sky130_fd_sc_hd__o211ai_4 _28404_ (.A1(net452),
    .A2(_06070_),
    .B1(_06072_),
    .C1(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__buf_6 _28405_ (.A(_05586_),
    .X(_06076_));
 sky130_fd_sc_hd__buf_6 _28406_ (.A(_05842_),
    .X(_06077_));
 sky130_fd_sc_hd__a22oi_4 _28407_ (.A1(_06076_),
    .A2(_05493_),
    .B1(_06077_),
    .B2(_05548_),
    .Y(_06078_));
 sky130_fd_sc_hd__nor2_8 _28408_ (.A(_05551_),
    .B(_06070_),
    .Y(_06079_));
 sky130_fd_sc_hd__o21ai_2 _28409_ (.A1(_06078_),
    .A2(_06079_),
    .B1(_06071_),
    .Y(_06080_));
 sky130_fd_sc_hd__o211ai_4 _28410_ (.A1(_06026_),
    .A2(_06069_),
    .B1(_06075_),
    .C1(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__o21a_1 _28411_ (.A1(_06023_),
    .A2(_06025_),
    .B1(_06016_),
    .X(_06082_));
 sky130_fd_sc_hd__o211ai_4 _28412_ (.A1(net452),
    .A2(_06070_),
    .B1(_06071_),
    .C1(_06074_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_2 _28413_ (.A1(_06078_),
    .A2(_06079_),
    .B1(_06072_),
    .Y(_06084_));
 sky130_fd_sc_hd__o211ai_4 _28414_ (.A1(_06021_),
    .A2(_06082_),
    .B1(_06083_),
    .C1(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__nor2_4 _28415_ (.A(_05932_),
    .B(_05929_),
    .Y(_06086_));
 sky130_fd_sc_hd__o2bb2ai_4 _28416_ (.A1_N(_06081_),
    .A2_N(_06085_),
    .B1(_05935_),
    .B2(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__nor2_2 _28417_ (.A(_05935_),
    .B(_06086_),
    .Y(_06088_));
 sky130_fd_sc_hd__nand3_4 _28418_ (.A(_06081_),
    .B(_06085_),
    .C(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__a21oi_4 _28419_ (.A1(_06087_),
    .A2(_06089_),
    .B1(_06035_),
    .Y(_06090_));
 sky130_fd_sc_hd__and3_1 _28420_ (.A(_06087_),
    .B(_06035_),
    .C(_06089_),
    .X(_06091_));
 sky130_fd_sc_hd__a21boi_4 _28421_ (.A1(_05940_),
    .A2(_05941_),
    .B1_N(_05937_),
    .Y(_06092_));
 sky130_fd_sc_hd__o21ai_4 _28422_ (.A1(_06090_),
    .A2(_06091_),
    .B1(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__a21o_1 _28423_ (.A1(_06087_),
    .A2(_06089_),
    .B1(_06035_),
    .X(_06094_));
 sky130_vsdinv _28424_ (.A(_06092_),
    .Y(_06095_));
 sky130_fd_sc_hd__nand3_4 _28425_ (.A(_06087_),
    .B(_06035_),
    .C(_06089_),
    .Y(_06096_));
 sky130_fd_sc_hd__nand3_4 _28426_ (.A(_06094_),
    .B(_06095_),
    .C(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__a21oi_4 _28427_ (.A1(_06093_),
    .A2(_06097_),
    .B1(_05953_),
    .Y(_06098_));
 sky130_fd_sc_hd__and3_2 _28428_ (.A(_06093_),
    .B(_05953_),
    .C(_06097_),
    .X(_06099_));
 sky130_fd_sc_hd__a22oi_4 _28429_ (.A1(_19671_),
    .A2(_05808_),
    .B1(_05780_),
    .B2(_19905_),
    .Y(_06100_));
 sky130_fd_sc_hd__nand3_4 _28430_ (.A(_05778_),
    .B(_05169_),
    .C(_19907_),
    .Y(_06101_));
 sky130_fd_sc_hd__nor2_8 _28431_ (.A(net447),
    .B(_06101_),
    .Y(_06102_));
 sky130_fd_sc_hd__nand2_4 _28432_ (.A(net476),
    .B(_19891_),
    .Y(_06103_));
 sky130_fd_sc_hd__o21ai_2 _28433_ (.A1(_06100_),
    .A2(_06102_),
    .B1(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__buf_4 _28434_ (.A(_05463_),
    .X(_06105_));
 sky130_fd_sc_hd__buf_6 _28435_ (.A(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__a22o_2 _28436_ (.A1(_05791_),
    .A2(_06106_),
    .B1(_05780_),
    .B2(_19905_),
    .X(_06107_));
 sky130_vsdinv _28437_ (.A(_06103_),
    .Y(_06108_));
 sky130_fd_sc_hd__nand3b_2 _28438_ (.A_N(_06102_),
    .B(_06107_),
    .C(_06108_),
    .Y(_06109_));
 sky130_fd_sc_hd__o2111ai_4 _28439_ (.A1(_05966_),
    .A2(_05960_),
    .B1(_05967_),
    .C1(_06104_),
    .D1(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__o21ai_2 _28440_ (.A1(_06100_),
    .A2(_06102_),
    .B1(_06108_),
    .Y(_06111_));
 sky130_fd_sc_hd__o21ai_2 _28441_ (.A1(_05966_),
    .A2(_05960_),
    .B1(_05967_),
    .Y(_06112_));
 sky130_fd_sc_hd__o211ai_4 _28442_ (.A1(_05981_),
    .A2(_06101_),
    .B1(_06103_),
    .C1(_06107_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand3_4 _28443_ (.A(_06111_),
    .B(_06112_),
    .C(_06113_),
    .Y(_06114_));
 sky130_fd_sc_hd__clkbuf_4 _28444_ (.A(\pcpi_mul.rs1[12] ),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_8 _28445_ (.A(_06115_),
    .X(_06116_));
 sky130_fd_sc_hd__clkbuf_2 _28446_ (.A(\pcpi_mul.rs1[11] ),
    .X(_06117_));
 sky130_fd_sc_hd__buf_4 _28447_ (.A(_06117_),
    .X(_06118_));
 sky130_fd_sc_hd__buf_6 _28448_ (.A(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__and4_4 _28449_ (.A(_05117_),
    .B(_05239_),
    .C(_06116_),
    .D(_06119_),
    .X(_06120_));
 sky130_fd_sc_hd__nand2_2 _28450_ (.A(_05157_),
    .B(_19902_),
    .Y(_06121_));
 sky130_fd_sc_hd__a22o_1 _28451_ (.A1(_05162_),
    .A2(_19899_),
    .B1(_05164_),
    .B2(_19895_),
    .X(_06122_));
 sky130_fd_sc_hd__nand3b_2 _28452_ (.A_N(_06120_),
    .B(_06121_),
    .C(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__a22oi_4 _28453_ (.A1(_05162_),
    .A2(_19899_),
    .B1(_05164_),
    .B2(_19895_),
    .Y(_06124_));
 sky130_vsdinv _28454_ (.A(_06121_),
    .Y(_06125_));
 sky130_fd_sc_hd__o21ai_2 _28455_ (.A1(_06124_),
    .A2(_06120_),
    .B1(_06125_),
    .Y(_06126_));
 sky130_fd_sc_hd__nand2_4 _28456_ (.A(_06123_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__a21o_1 _28457_ (.A1(_06110_),
    .A2(_06114_),
    .B1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__nand3_4 _28458_ (.A(_06110_),
    .B(_06114_),
    .C(_06127_),
    .Y(_06129_));
 sky130_fd_sc_hd__nand2_1 _28459_ (.A(_06128_),
    .B(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__a21oi_2 _28460_ (.A1(_05964_),
    .A2(_05968_),
    .B1(_05969_),
    .Y(_06131_));
 sky130_fd_sc_hd__o21a_1 _28461_ (.A1(_05988_),
    .A2(_06131_),
    .B1(_05970_),
    .X(_06132_));
 sky130_vsdinv _28462_ (.A(_05985_),
    .Y(_06133_));
 sky130_fd_sc_hd__nor2_2 _28463_ (.A(_05978_),
    .B(_06133_),
    .Y(_06134_));
 sky130_fd_sc_hd__a21oi_2 _28464_ (.A1(_06130_),
    .A2(_06132_),
    .B1(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__o21ai_2 _28465_ (.A1(_05988_),
    .A2(_06131_),
    .B1(_05970_),
    .Y(_06136_));
 sky130_fd_sc_hd__nand3_4 _28466_ (.A(_06136_),
    .B(_06128_),
    .C(_06129_),
    .Y(_06137_));
 sky130_fd_sc_hd__a21oi_2 _28467_ (.A1(_06110_),
    .A2(_06114_),
    .B1(_06127_),
    .Y(_06138_));
 sky130_fd_sc_hd__and3_1 _28468_ (.A(_06110_),
    .B(_06114_),
    .C(_06127_),
    .X(_06139_));
 sky130_fd_sc_hd__o21ai_4 _28469_ (.A1(_06138_),
    .A2(_06139_),
    .B1(_06132_),
    .Y(_06140_));
 sky130_vsdinv _28470_ (.A(_06134_),
    .Y(_06141_));
 sky130_fd_sc_hd__a21oi_2 _28471_ (.A1(_06140_),
    .A2(_06137_),
    .B1(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__a21oi_4 _28472_ (.A1(_06135_),
    .A2(_06137_),
    .B1(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__o21ai_2 _28473_ (.A1(_06098_),
    .A2(_06099_),
    .B1(_06143_),
    .Y(_06144_));
 sky130_fd_sc_hd__o2bb2ai_4 _28474_ (.A1_N(_06097_),
    .A2_N(_06093_),
    .B1(_05944_),
    .B2(_05947_),
    .Y(_06145_));
 sky130_fd_sc_hd__nand3_2 _28475_ (.A(_06093_),
    .B(_05953_),
    .C(_06097_),
    .Y(_06146_));
 sky130_fd_sc_hd__a21o_1 _28476_ (.A1(_06140_),
    .A2(_06137_),
    .B1(_06141_),
    .X(_06147_));
 sky130_fd_sc_hd__nand3_4 _28477_ (.A(_06140_),
    .B(_06141_),
    .C(_06137_),
    .Y(_06148_));
 sky130_fd_sc_hd__nand2_4 _28478_ (.A(_06147_),
    .B(_06148_),
    .Y(_06149_));
 sky130_fd_sc_hd__nand3_2 _28479_ (.A(_06145_),
    .B(_06146_),
    .C(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__nand3b_4 _28480_ (.A_N(_06068_),
    .B(_06144_),
    .C(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__o21ai_2 _28481_ (.A1(_06098_),
    .A2(_06099_),
    .B1(_06149_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand3_2 _28482_ (.A(_06145_),
    .B(_06143_),
    .C(_06146_),
    .Y(_06153_));
 sky130_fd_sc_hd__nand3_4 _28483_ (.A(_06152_),
    .B(_06153_),
    .C(_06068_),
    .Y(_06154_));
 sky130_fd_sc_hd__nand2_2 _28484_ (.A(_06151_),
    .B(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__buf_6 _28485_ (.A(_19651_),
    .X(_06156_));
 sky130_fd_sc_hd__nand2_2 _28486_ (.A(_06156_),
    .B(_05230_),
    .Y(_06157_));
 sky130_fd_sc_hd__clkbuf_4 _28487_ (.A(\pcpi_mul.rs2[10] ),
    .X(_06158_));
 sky130_fd_sc_hd__buf_6 _28488_ (.A(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_8 _28489_ (.A(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__nand3b_4 _28490_ (.A_N(_06157_),
    .B(_06160_),
    .C(_19925_),
    .Y(_06161_));
 sky130_fd_sc_hd__nand2_1 _28491_ (.A(_19655_),
    .B(_05147_),
    .Y(_06162_));
 sky130_fd_sc_hd__nand2_2 _28492_ (.A(_06157_),
    .B(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__nand2_2 _28493_ (.A(_06014_),
    .B(_05237_),
    .Y(_06164_));
 sky130_fd_sc_hd__a21o_1 _28494_ (.A1(_06161_),
    .A2(_06163_),
    .B1(_06164_),
    .X(_06165_));
 sky130_fd_sc_hd__nand3_4 _28495_ (.A(_06161_),
    .B(_06163_),
    .C(_06164_),
    .Y(_06166_));
 sky130_fd_sc_hd__clkbuf_4 _28496_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06167_));
 sky130_fd_sc_hd__buf_2 _28497_ (.A(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__buf_8 _28498_ (.A(_06168_),
    .X(_06169_));
 sky130_fd_sc_hd__nand2_1 _28499_ (.A(_06169_),
    .B(_05213_),
    .Y(_06170_));
 sky130_fd_sc_hd__nand2_1 _28500_ (.A(_19650_),
    .B(_05123_),
    .Y(_06171_));
 sky130_fd_sc_hd__or2_2 _28501_ (.A(_06170_),
    .B(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__nand2_1 _28502_ (.A(_06170_),
    .B(_06171_),
    .Y(_06173_));
 sky130_fd_sc_hd__nand2_2 _28503_ (.A(_06172_),
    .B(_06173_),
    .Y(_06174_));
 sky130_fd_sc_hd__a21oi_4 _28504_ (.A1(_06165_),
    .A2(_06166_),
    .B1(_06174_),
    .Y(_06175_));
 sky130_fd_sc_hd__and3_1 _28505_ (.A(_06165_),
    .B(_06174_),
    .C(_06166_),
    .X(_06176_));
 sky130_fd_sc_hd__or2_4 _28506_ (.A(_06175_),
    .B(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__nand2_2 _28507_ (.A(_06155_),
    .B(_06177_),
    .Y(_06178_));
 sky130_vsdinv _28508_ (.A(_06177_),
    .Y(_06179_));
 sky130_fd_sc_hd__nand3_4 _28509_ (.A(_06151_),
    .B(_06154_),
    .C(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__nand2_1 _28510_ (.A(_06178_),
    .B(_06180_),
    .Y(_06181_));
 sky130_fd_sc_hd__nand2_1 _28511_ (.A(_06181_),
    .B(_06038_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand3b_4 _28512_ (.A_N(_06038_),
    .B(_06178_),
    .C(_06180_),
    .Y(_06183_));
 sky130_fd_sc_hd__nand2_1 _28513_ (.A(_06182_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__and2_1 _28514_ (.A(_05998_),
    .B(_05993_),
    .X(_06185_));
 sky130_fd_sc_hd__nor2_4 _28515_ (.A(_06185_),
    .B(_06006_),
    .Y(_06186_));
 sky130_fd_sc_hd__and2_1 _28516_ (.A(_06006_),
    .B(_06185_),
    .X(_06187_));
 sky130_fd_sc_hd__or2_1 _28517_ (.A(_06186_),
    .B(_06187_),
    .X(_06188_));
 sky130_vsdinv _28518_ (.A(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_1 _28519_ (.A(_06184_),
    .B(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__a21oi_2 _28520_ (.A1(_06049_),
    .A2(_06045_),
    .B1(_06040_),
    .Y(_06191_));
 sky130_fd_sc_hd__nand3_1 _28521_ (.A(_06182_),
    .B(_06188_),
    .C(_06183_),
    .Y(_06192_));
 sky130_fd_sc_hd__nand3_2 _28522_ (.A(_06190_),
    .B(_06191_),
    .C(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__and2_1 _28523_ (.A(_06193_),
    .B(_06043_),
    .X(_06194_));
 sky130_vsdinv _28524_ (.A(_06183_),
    .Y(_06195_));
 sky130_fd_sc_hd__nand2_1 _28525_ (.A(_06182_),
    .B(_06189_),
    .Y(_06196_));
 sky130_vsdinv _28526_ (.A(_06191_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_1 _28527_ (.A(_06184_),
    .B(_06188_),
    .Y(_06198_));
 sky130_fd_sc_hd__o211ai_2 _28528_ (.A1(_06195_),
    .A2(_06196_),
    .B1(_06197_),
    .C1(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__a21oi_1 _28529_ (.A1(_06199_),
    .A2(_06193_),
    .B1(_06043_),
    .Y(_06200_));
 sky130_fd_sc_hd__nand2_1 _28530_ (.A(_06054_),
    .B(_06058_),
    .Y(_06201_));
 sky130_fd_sc_hd__o21bai_1 _28531_ (.A1(_06194_),
    .A2(_06200_),
    .B1_N(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__a21o_1 _28532_ (.A1(_06199_),
    .A2(_06193_),
    .B1(_06043_),
    .X(_06203_));
 sky130_fd_sc_hd__nand2_1 _28533_ (.A(_06193_),
    .B(_06043_),
    .Y(_06204_));
 sky130_fd_sc_hd__nand3_1 _28534_ (.A(_06203_),
    .B(_06201_),
    .C(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__nand2_1 _28535_ (.A(_06202_),
    .B(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__a22oi_4 _28536_ (.A1(_06054_),
    .A2(_06062_),
    .B1(_06067_),
    .B2(_06065_),
    .Y(_06207_));
 sky130_fd_sc_hd__xor2_1 _28537_ (.A(_06206_),
    .B(_06207_),
    .X(_02632_));
 sky130_fd_sc_hd__nand2_1 _28538_ (.A(_06196_),
    .B(_06183_),
    .Y(_06208_));
 sky130_fd_sc_hd__and2_2 _28539_ (.A(_06148_),
    .B(_06137_),
    .X(_06209_));
 sky130_fd_sc_hd__nor2_8 _28540_ (.A(_06209_),
    .B(_06154_),
    .Y(_06210_));
 sky130_fd_sc_hd__and2_2 _28541_ (.A(_06154_),
    .B(_06209_),
    .X(_06211_));
 sky130_fd_sc_hd__nor2_8 _28542_ (.A(_06210_),
    .B(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__a22oi_4 _28543_ (.A1(_05837_),
    .A2(_05548_),
    .B1(_06077_),
    .B2(_05666_),
    .Y(_06213_));
 sky130_vsdinv _28544_ (.A(\pcpi_mul.rs1[7] ),
    .Y(_06214_));
 sky130_fd_sc_hd__buf_4 _28545_ (.A(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__buf_4 _28546_ (.A(\pcpi_mul.rs2[7] ),
    .X(_06216_));
 sky130_fd_sc_hd__buf_4 _28547_ (.A(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__nand3_4 _28548_ (.A(_05451_),
    .B(_06217_),
    .C(_05656_),
    .Y(_06218_));
 sky130_fd_sc_hd__nor2_8 _28549_ (.A(net472),
    .B(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__nand2_2 _28550_ (.A(_05835_),
    .B(_05958_),
    .Y(_06220_));
 sky130_fd_sc_hd__o21ai_2 _28551_ (.A1(_06213_),
    .A2(_06219_),
    .B1(_06220_),
    .Y(_06221_));
 sky130_vsdinv _28552_ (.A(_06220_),
    .Y(_06222_));
 sky130_fd_sc_hd__a22o_2 _28553_ (.A1(_05841_),
    .A2(_19914_),
    .B1(_05843_),
    .B2(_05671_),
    .X(_06223_));
 sky130_fd_sc_hd__o211ai_4 _28554_ (.A1(net472),
    .A2(_06218_),
    .B1(_06222_),
    .C1(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__a22oi_4 _28555_ (.A1(_19653_),
    .A2(_19928_),
    .B1(net457),
    .B2(_19925_),
    .Y(_06225_));
 sky130_fd_sc_hd__o21ai_2 _28556_ (.A1(_06164_),
    .A2(_06225_),
    .B1(_06161_),
    .Y(_06226_));
 sky130_fd_sc_hd__nand3_4 _28557_ (.A(_06221_),
    .B(_06224_),
    .C(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__o21ai_2 _28558_ (.A1(_06213_),
    .A2(_06219_),
    .B1(_06222_),
    .Y(_06228_));
 sky130_fd_sc_hd__o21ai_1 _28559_ (.A1(_06157_),
    .A2(_06162_),
    .B1(_06164_),
    .Y(_06229_));
 sky130_fd_sc_hd__nand2_1 _28560_ (.A(_06229_),
    .B(_06163_),
    .Y(_06230_));
 sky130_fd_sc_hd__o211ai_2 _28561_ (.A1(net472),
    .A2(_06218_),
    .B1(_06220_),
    .C1(_06223_),
    .Y(_06231_));
 sky130_fd_sc_hd__nand3_4 _28562_ (.A(_06228_),
    .B(_06230_),
    .C(_06231_),
    .Y(_06232_));
 sky130_fd_sc_hd__nor2_8 _28563_ (.A(_06072_),
    .B(_06079_),
    .Y(_06233_));
 sky130_fd_sc_hd__o2bb2ai_4 _28564_ (.A1_N(_06227_),
    .A2_N(_06232_),
    .B1(_06078_),
    .B2(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__nor2_2 _28565_ (.A(_06078_),
    .B(_06233_),
    .Y(_06235_));
 sky130_fd_sc_hd__nand3_4 _28566_ (.A(_06227_),
    .B(_06232_),
    .C(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__a21oi_4 _28567_ (.A1(_06234_),
    .A2(_06236_),
    .B1(_06175_),
    .Y(_06237_));
 sky130_fd_sc_hd__and3_1 _28568_ (.A(_06221_),
    .B(_06226_),
    .C(_06224_),
    .X(_06238_));
 sky130_fd_sc_hd__nand2_1 _28569_ (.A(_06232_),
    .B(_06235_),
    .Y(_06239_));
 sky130_fd_sc_hd__o211a_1 _28570_ (.A1(_06238_),
    .A2(_06239_),
    .B1(_06175_),
    .C1(_06234_),
    .X(_06240_));
 sky130_vsdinv _28571_ (.A(_06081_),
    .Y(_06241_));
 sky130_fd_sc_hd__a21oi_1 _28572_ (.A1(_06085_),
    .A2(_06088_),
    .B1(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__buf_2 _28573_ (.A(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__o21ai_2 _28574_ (.A1(_06237_),
    .A2(_06240_),
    .B1(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__o21ai_2 _28575_ (.A1(_06092_),
    .A2(_06090_),
    .B1(_06096_),
    .Y(_06245_));
 sky130_fd_sc_hd__nand2_1 _28576_ (.A(_06234_),
    .B(_06236_),
    .Y(_06246_));
 sky130_vsdinv _28577_ (.A(_06175_),
    .Y(_06247_));
 sky130_fd_sc_hd__nand2_2 _28578_ (.A(_06246_),
    .B(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__nand3_4 _28579_ (.A(_06234_),
    .B(_06175_),
    .C(_06236_),
    .Y(_06249_));
 sky130_fd_sc_hd__nand3b_4 _28580_ (.A_N(_06243_),
    .B(_06248_),
    .C(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__nand3_4 _28581_ (.A(_06244_),
    .B(_06245_),
    .C(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__o21bai_2 _28582_ (.A1(_06237_),
    .A2(_06240_),
    .B1_N(_06242_),
    .Y(_06252_));
 sky130_fd_sc_hd__nand2_1 _28583_ (.A(_06096_),
    .B(_06092_),
    .Y(_06253_));
 sky130_fd_sc_hd__nand2_1 _28584_ (.A(_06253_),
    .B(_06094_),
    .Y(_06254_));
 sky130_fd_sc_hd__nand3_2 _28585_ (.A(_06248_),
    .B(_06249_),
    .C(_06243_),
    .Y(_06255_));
 sky130_fd_sc_hd__nand3_4 _28586_ (.A(_06252_),
    .B(_06254_),
    .C(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__buf_6 _28587_ (.A(_05558_),
    .X(_06257_));
 sky130_fd_sc_hd__buf_6 _28588_ (.A(_19672_),
    .X(_06258_));
 sky130_fd_sc_hd__buf_4 _28589_ (.A(_05642_),
    .X(_06259_));
 sky130_fd_sc_hd__buf_4 _28590_ (.A(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__a22oi_4 _28591_ (.A1(_05778_),
    .A2(_06257_),
    .B1(_06258_),
    .B2(_06260_),
    .Y(_06261_));
 sky130_vsdinv _28592_ (.A(_05642_),
    .Y(_06262_));
 sky130_fd_sc_hd__buf_2 _28593_ (.A(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__buf_4 _28594_ (.A(_19903_),
    .X(_06264_));
 sky130_fd_sc_hd__nand3_4 _28595_ (.A(_05203_),
    .B(_05285_),
    .C(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__nor2_8 _28596_ (.A(_06263_),
    .B(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__buf_6 _28597_ (.A(_19886_),
    .X(_06267_));
 sky130_fd_sc_hd__nand2_4 _28598_ (.A(net495),
    .B(_06267_),
    .Y(_06268_));
 sky130_vsdinv _28599_ (.A(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__o21ai_4 _28600_ (.A1(_06261_),
    .A2(_06266_),
    .B1(_06269_),
    .Y(_06270_));
 sky130_fd_sc_hd__a21oi_4 _28601_ (.A1(_06107_),
    .A2(_06108_),
    .B1(_06102_),
    .Y(_06271_));
 sky130_fd_sc_hd__buf_6 _28602_ (.A(_06263_),
    .X(_06272_));
 sky130_fd_sc_hd__a22o_2 _28603_ (.A1(_05778_),
    .A2(_06257_),
    .B1(_19673_),
    .B2(_06260_),
    .X(_06273_));
 sky130_fd_sc_hd__o211ai_4 _28604_ (.A1(_06272_),
    .A2(_06265_),
    .B1(_06268_),
    .C1(_06273_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand3_4 _28605_ (.A(_06270_),
    .B(_06271_),
    .C(_06274_),
    .Y(_06275_));
 sky130_fd_sc_hd__nor2_2 _28606_ (.A(_06103_),
    .B(_06100_),
    .Y(_06276_));
 sky130_fd_sc_hd__o211ai_4 _28607_ (.A1(_06272_),
    .A2(_06265_),
    .B1(_06269_),
    .C1(_06273_),
    .Y(_06277_));
 sky130_fd_sc_hd__o21ai_2 _28608_ (.A1(_06261_),
    .A2(_06266_),
    .B1(_06268_),
    .Y(_06278_));
 sky130_fd_sc_hd__o211ai_4 _28609_ (.A1(_06102_),
    .A2(_06276_),
    .B1(_06277_),
    .C1(_06278_),
    .Y(_06279_));
 sky130_fd_sc_hd__nand2_4 _28610_ (.A(_05807_),
    .B(_19899_),
    .Y(_06280_));
 sky130_fd_sc_hd__buf_6 _28611_ (.A(_05161_),
    .X(_06281_));
 sky130_fd_sc_hd__clkbuf_4 _28612_ (.A(\pcpi_mul.rs1[13] ),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_4 _28613_ (.A(_06282_),
    .X(_06283_));
 sky130_fd_sc_hd__buf_6 _28614_ (.A(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__a22oi_4 _28615_ (.A1(_06281_),
    .A2(_19895_),
    .B1(_05235_),
    .B2(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__buf_6 _28616_ (.A(_06283_),
    .X(_06286_));
 sky130_fd_sc_hd__buf_2 _28617_ (.A(\pcpi_mul.rs1[12] ),
    .X(_06287_));
 sky130_fd_sc_hd__buf_4 _28618_ (.A(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__buf_6 _28619_ (.A(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__and4_4 _28620_ (.A(_06281_),
    .B(_05223_),
    .C(_06286_),
    .D(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__nor3_4 _28621_ (.A(_06280_),
    .B(_06285_),
    .C(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__o21a_1 _28622_ (.A1(_06285_),
    .A2(_06290_),
    .B1(_06280_),
    .X(_06292_));
 sky130_fd_sc_hd__o2bb2ai_2 _28623_ (.A1_N(_06275_),
    .A2_N(_06279_),
    .B1(_06291_),
    .B2(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__nor2_1 _28624_ (.A(_06285_),
    .B(_06290_),
    .Y(_06294_));
 sky130_fd_sc_hd__nand2_2 _28625_ (.A(_06294_),
    .B(_06280_),
    .Y(_06295_));
 sky130_fd_sc_hd__o21bai_2 _28626_ (.A1(_06285_),
    .A2(_06290_),
    .B1_N(_06280_),
    .Y(_06296_));
 sky130_fd_sc_hd__nand2_1 _28627_ (.A(_06295_),
    .B(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__nand3_2 _28628_ (.A(_06297_),
    .B(_06279_),
    .C(_06275_),
    .Y(_06298_));
 sky130_fd_sc_hd__nand2_1 _28629_ (.A(_06127_),
    .B(_06114_),
    .Y(_06299_));
 sky130_fd_sc_hd__nand2_2 _28630_ (.A(_06299_),
    .B(_06110_),
    .Y(_06300_));
 sky130_fd_sc_hd__a21oi_1 _28631_ (.A1(_06293_),
    .A2(_06298_),
    .B1(_06300_),
    .Y(_06301_));
 sky130_vsdinv _28632_ (.A(_06279_),
    .Y(_06302_));
 sky130_fd_sc_hd__nand2_2 _28633_ (.A(_06297_),
    .B(_06275_),
    .Y(_06303_));
 sky130_fd_sc_hd__o211a_1 _28634_ (.A1(_06302_),
    .A2(_06303_),
    .B1(_06293_),
    .C1(_06300_),
    .X(_06304_));
 sky130_fd_sc_hd__nor3_4 _28635_ (.A(_06121_),
    .B(_06124_),
    .C(_06120_),
    .Y(_06305_));
 sky130_fd_sc_hd__nor2_4 _28636_ (.A(_06120_),
    .B(_06305_),
    .Y(_06306_));
 sky130_vsdinv _28637_ (.A(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__o21ai_1 _28638_ (.A1(_06301_),
    .A2(_06304_),
    .B1(_06307_),
    .Y(_06308_));
 sky130_fd_sc_hd__a21o_1 _28639_ (.A1(_06293_),
    .A2(_06298_),
    .B1(_06300_),
    .X(_06309_));
 sky130_fd_sc_hd__nand3_2 _28640_ (.A(_06300_),
    .B(_06293_),
    .C(_06298_),
    .Y(_06310_));
 sky130_fd_sc_hd__nand3_1 _28641_ (.A(_06309_),
    .B(_06306_),
    .C(_06310_),
    .Y(_06311_));
 sky130_fd_sc_hd__nand2_2 _28642_ (.A(_06308_),
    .B(_06311_),
    .Y(_06312_));
 sky130_fd_sc_hd__a21oi_1 _28643_ (.A1(_06251_),
    .A2(_06256_),
    .B1(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__a21oi_1 _28644_ (.A1(_06309_),
    .A2(_06310_),
    .B1(_06306_),
    .Y(_06314_));
 sky130_fd_sc_hd__and3_1 _28645_ (.A(_06309_),
    .B(_06306_),
    .C(_06310_),
    .X(_06315_));
 sky130_fd_sc_hd__o211a_1 _28646_ (.A1(_06314_),
    .A2(_06315_),
    .B1(_06256_),
    .C1(_06251_),
    .X(_06316_));
 sky130_fd_sc_hd__a21oi_4 _28647_ (.A1(_06145_),
    .A2(_06143_),
    .B1(_06099_),
    .Y(_06317_));
 sky130_fd_sc_hd__o21ai_2 _28648_ (.A1(_06313_),
    .A2(_06316_),
    .B1(_06317_),
    .Y(_06318_));
 sky130_vsdinv _28649_ (.A(_06097_),
    .Y(_06319_));
 sky130_fd_sc_hd__nand2_1 _28650_ (.A(_06093_),
    .B(_05953_),
    .Y(_06320_));
 sky130_fd_sc_hd__o22ai_4 _28651_ (.A1(_06319_),
    .A2(_06320_),
    .B1(_06149_),
    .B2(_06098_),
    .Y(_06321_));
 sky130_fd_sc_hd__nand3_4 _28652_ (.A(_06312_),
    .B(_06251_),
    .C(_06256_),
    .Y(_06322_));
 sky130_fd_sc_hd__a21o_1 _28653_ (.A1(_06251_),
    .A2(_06256_),
    .B1(_06312_),
    .X(_06323_));
 sky130_fd_sc_hd__nand3_4 _28654_ (.A(_06321_),
    .B(_06322_),
    .C(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__buf_6 _28655_ (.A(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__buf_4 _28656_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06326_));
 sky130_fd_sc_hd__clkbuf_8 _28657_ (.A(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__a22oi_4 _28658_ (.A1(_06327_),
    .A2(_06015_),
    .B1(net448),
    .B2(_05237_),
    .Y(_06328_));
 sky130_fd_sc_hd__nand2_2 _28659_ (.A(_06022_),
    .B(_05359_),
    .Y(_06329_));
 sky130_fd_sc_hd__buf_6 _28660_ (.A(_05272_),
    .X(_06330_));
 sky130_fd_sc_hd__nand2_1 _28661_ (.A(_06159_),
    .B(_06330_),
    .Y(_06331_));
 sky130_fd_sc_hd__nor2_1 _28662_ (.A(_06329_),
    .B(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand2_2 _28663_ (.A(_06014_),
    .B(_06073_),
    .Y(_06333_));
 sky130_fd_sc_hd__o21bai_2 _28664_ (.A1(_06328_),
    .A2(_06332_),
    .B1_N(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__buf_6 _28665_ (.A(_05735_),
    .X(_06335_));
 sky130_fd_sc_hd__clkbuf_8 _28666_ (.A(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__nand3b_4 _28667_ (.A_N(_06329_),
    .B(_06336_),
    .C(_19921_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_1 _28668_ (.A(_06329_),
    .B(_06331_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand3_2 _28669_ (.A(_06337_),
    .B(_06333_),
    .C(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__nand2_4 _28670_ (.A(_06334_),
    .B(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__buf_6 _28671_ (.A(_19643_),
    .X(_06341_));
 sky130_fd_sc_hd__buf_6 _28672_ (.A(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__clkbuf_8 _28673_ (.A(_06168_),
    .X(_06343_));
 sky130_fd_sc_hd__a22oi_4 _28674_ (.A1(_06342_),
    .A2(_05406_),
    .B1(_06343_),
    .B2(_05158_),
    .Y(_06344_));
 sky130_fd_sc_hd__buf_6 _28675_ (.A(_06167_),
    .X(_06345_));
 sky130_fd_sc_hd__nand2_2 _28676_ (.A(_06345_),
    .B(_19930_),
    .Y(_06346_));
 sky130_fd_sc_hd__nand2_2 _28677_ (.A(_19644_),
    .B(_19933_),
    .Y(_06347_));
 sky130_fd_sc_hd__nor2_2 _28678_ (.A(_06346_),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__buf_6 _28679_ (.A(_19649_),
    .X(_06349_));
 sky130_fd_sc_hd__nand2_2 _28680_ (.A(_06349_),
    .B(_05121_),
    .Y(_06350_));
 sky130_fd_sc_hd__o21ai_2 _28681_ (.A1(_06344_),
    .A2(_06348_),
    .B1(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__clkbuf_2 _28682_ (.A(_19644_),
    .X(_06352_));
 sky130_fd_sc_hd__nand3b_4 _28683_ (.A_N(_06346_),
    .B(_06352_),
    .C(_05406_),
    .Y(_06353_));
 sky130_vsdinv _28684_ (.A(_06350_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand2_2 _28685_ (.A(_06346_),
    .B(_06347_),
    .Y(_06355_));
 sky130_fd_sc_hd__nand3_2 _28686_ (.A(_06353_),
    .B(_06354_),
    .C(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__nand3b_4 _28687_ (.A_N(_06172_),
    .B(_06351_),
    .C(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__o21ai_2 _28688_ (.A1(_06344_),
    .A2(_06348_),
    .B1(_06354_),
    .Y(_06358_));
 sky130_fd_sc_hd__nand3_2 _28689_ (.A(_06353_),
    .B(_06350_),
    .C(_06355_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand3_4 _28690_ (.A(_06358_),
    .B(_06359_),
    .C(_06172_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand2_1 _28691_ (.A(_06357_),
    .B(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__nor2_1 _28692_ (.A(_06340_),
    .B(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__and2_1 _28693_ (.A(_06361_),
    .B(_06340_),
    .X(_06363_));
 sky130_fd_sc_hd__or2_2 _28694_ (.A(_06362_),
    .B(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__a21oi_4 _28695_ (.A1(_06318_),
    .A2(_06325_),
    .B1(_06364_),
    .Y(_06365_));
 sky130_fd_sc_hd__nor2_4 _28696_ (.A(_06180_),
    .B(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__nand2_1 _28697_ (.A(_06323_),
    .B(_06322_),
    .Y(_06367_));
 sky130_vsdinv _28698_ (.A(_06364_),
    .Y(_06368_));
 sky130_fd_sc_hd__a21oi_4 _28699_ (.A1(_06367_),
    .A2(_06317_),
    .B1(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__nand2_2 _28700_ (.A(_06369_),
    .B(_06325_),
    .Y(_06370_));
 sky130_fd_sc_hd__nand2_1 _28701_ (.A(_06366_),
    .B(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__o211a_2 _28702_ (.A1(_06362_),
    .A2(_06363_),
    .B1(_06325_),
    .C1(_06318_),
    .X(_06372_));
 sky130_fd_sc_hd__o22ai_4 _28703_ (.A1(_06177_),
    .A2(_06155_),
    .B1(_06365_),
    .B2(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__nand2_1 _28704_ (.A(_06371_),
    .B(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__nor2_2 _28705_ (.A(_06212_),
    .B(_06374_),
    .Y(_06375_));
 sky130_vsdinv _28706_ (.A(_06375_),
    .Y(_06376_));
 sky130_fd_sc_hd__nand2_1 _28707_ (.A(_06374_),
    .B(_06212_),
    .Y(_06377_));
 sky130_fd_sc_hd__nand3b_2 _28708_ (.A_N(_06208_),
    .B(_06376_),
    .C(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_2 _28709_ (.A(_06378_),
    .B(_06186_),
    .Y(_06379_));
 sky130_vsdinv _28710_ (.A(_06377_),
    .Y(_06380_));
 sky130_fd_sc_hd__o21ai_2 _28711_ (.A1(_06375_),
    .A2(_06380_),
    .B1(_06208_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2_1 _28712_ (.A(_06381_),
    .B(_06378_),
    .Y(_06382_));
 sky130_vsdinv _28713_ (.A(_06186_),
    .Y(_06383_));
 sky130_fd_sc_hd__nand2_1 _28714_ (.A(_06204_),
    .B(_06199_),
    .Y(_06384_));
 sky130_fd_sc_hd__a21boi_2 _28715_ (.A1(_06382_),
    .A2(_06383_),
    .B1_N(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__nand2_1 _28716_ (.A(_06382_),
    .B(_06383_),
    .Y(_06386_));
 sky130_fd_sc_hd__a21oi_1 _28717_ (.A1(_06386_),
    .A2(_06379_),
    .B1(_06384_),
    .Y(_06387_));
 sky130_fd_sc_hd__a21oi_2 _28718_ (.A1(_06379_),
    .A2(_06385_),
    .B1(_06387_),
    .Y(_06388_));
 sky130_vsdinv _28719_ (.A(_06205_),
    .Y(_06389_));
 sky130_fd_sc_hd__o21bai_1 _28720_ (.A1(_06206_),
    .A2(_06207_),
    .B1_N(_06389_),
    .Y(_06390_));
 sky130_fd_sc_hd__or2_1 _28721_ (.A(_06388_),
    .B(_06390_),
    .X(_06391_));
 sky130_fd_sc_hd__nand2_2 _28722_ (.A(_06390_),
    .B(_06388_),
    .Y(_06392_));
 sky130_fd_sc_hd__and2_1 _28723_ (.A(_06391_),
    .B(_06392_),
    .X(_02633_));
 sky130_fd_sc_hd__nand2_2 _28724_ (.A(_06379_),
    .B(_06381_),
    .Y(_06393_));
 sky130_fd_sc_hd__a21oi_4 _28725_ (.A1(_06309_),
    .A2(_06307_),
    .B1(_06304_),
    .Y(_06394_));
 sky130_vsdinv _28726_ (.A(_06394_),
    .Y(_06395_));
 sky130_fd_sc_hd__and2_4 _28727_ (.A(_06324_),
    .B(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__nor2_8 _28728_ (.A(_06395_),
    .B(_06325_),
    .Y(_06397_));
 sky130_fd_sc_hd__buf_6 _28729_ (.A(_19651_),
    .X(_06398_));
 sky130_fd_sc_hd__buf_6 _28730_ (.A(_19654_),
    .X(_06399_));
 sky130_fd_sc_hd__a22oi_4 _28731_ (.A1(_06398_),
    .A2(_05225_),
    .B1(_06399_),
    .B2(_06073_),
    .Y(_06400_));
 sky130_fd_sc_hd__buf_4 _28732_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06401_));
 sky130_fd_sc_hd__nand2_2 _28733_ (.A(_06401_),
    .B(_05224_),
    .Y(_06402_));
 sky130_fd_sc_hd__nand2_1 _28734_ (.A(_06335_),
    .B(_05378_),
    .Y(_06403_));
 sky130_fd_sc_hd__nor2_1 _28735_ (.A(_06402_),
    .B(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__nand2_2 _28736_ (.A(_19659_),
    .B(_05548_),
    .Y(_06405_));
 sky130_fd_sc_hd__o21bai_2 _28737_ (.A1(_06400_),
    .A2(_06404_),
    .B1_N(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand3b_4 _28738_ (.A_N(_06402_),
    .B(net448),
    .C(_19918_),
    .Y(_06407_));
 sky130_fd_sc_hd__nand2_1 _28739_ (.A(_06402_),
    .B(_06403_),
    .Y(_06408_));
 sky130_fd_sc_hd__nand3_2 _28740_ (.A(_06407_),
    .B(_06408_),
    .C(_06405_),
    .Y(_06409_));
 sky130_fd_sc_hd__nand2_4 _28741_ (.A(_06406_),
    .B(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__buf_8 _28742_ (.A(_06341_),
    .X(_06411_));
 sky130_fd_sc_hd__a22oi_4 _28743_ (.A1(_06411_),
    .A2(_05158_),
    .B1(_06343_),
    .B2(_05128_),
    .Y(_06412_));
 sky130_fd_sc_hd__clkbuf_4 _28744_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06413_));
 sky130_fd_sc_hd__buf_6 _28745_ (.A(_06413_),
    .X(_06414_));
 sky130_fd_sc_hd__nand2_2 _28746_ (.A(_06414_),
    .B(_05281_),
    .Y(_06415_));
 sky130_fd_sc_hd__buf_8 _28747_ (.A(_06167_),
    .X(_06416_));
 sky130_fd_sc_hd__nand2_2 _28748_ (.A(_06416_),
    .B(_06020_),
    .Y(_06417_));
 sky130_fd_sc_hd__nor2_1 _28749_ (.A(_06415_),
    .B(_06417_),
    .Y(_06418_));
 sky130_fd_sc_hd__buf_6 _28750_ (.A(\pcpi_mul.rs2[12] ),
    .X(_06419_));
 sky130_fd_sc_hd__nand2_2 _28751_ (.A(_06419_),
    .B(_05838_),
    .Y(_06420_));
 sky130_fd_sc_hd__o21bai_2 _28752_ (.A1(_06412_),
    .A2(_06418_),
    .B1_N(_06420_),
    .Y(_06421_));
 sky130_fd_sc_hd__clkbuf_8 _28753_ (.A(_19646_),
    .X(_06422_));
 sky130_fd_sc_hd__buf_8 _28754_ (.A(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__nand3b_2 _28755_ (.A_N(_06415_),
    .B(_06423_),
    .C(_19928_),
    .Y(_06424_));
 sky130_fd_sc_hd__nand2_2 _28756_ (.A(_06415_),
    .B(_06417_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand3_4 _28757_ (.A(_06424_),
    .B(_06425_),
    .C(_06420_),
    .Y(_06426_));
 sky130_fd_sc_hd__o21ai_1 _28758_ (.A1(_06346_),
    .A2(_06347_),
    .B1(_06350_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand2_2 _28759_ (.A(_06427_),
    .B(_06355_),
    .Y(_06428_));
 sky130_fd_sc_hd__a21o_1 _28760_ (.A1(_06421_),
    .A2(_06426_),
    .B1(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__nand3_2 _28761_ (.A(_06421_),
    .B(_06426_),
    .C(_06428_),
    .Y(_06430_));
 sky130_fd_sc_hd__nand2_2 _28762_ (.A(_06429_),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__xnor2_4 _28763_ (.A(_06410_),
    .B(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__inv_8 _28764_ (.A(_19640_),
    .Y(_06433_));
 sky130_fd_sc_hd__buf_2 _28765_ (.A(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__nor2_4 _28766_ (.A(_06434_),
    .B(_04842_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2_2 _28767_ (.A(_06432_),
    .B(_06435_),
    .Y(_06436_));
 sky130_vsdinv _28768_ (.A(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__nor2_4 _28769_ (.A(_06435_),
    .B(_06432_),
    .Y(_06438_));
 sky130_fd_sc_hd__a22oi_4 _28770_ (.A1(_05197_),
    .A2(_19901_),
    .B1(_05169_),
    .B2(_05774_),
    .Y(_06439_));
 sky130_fd_sc_hd__buf_4 _28771_ (.A(_06117_),
    .X(_06440_));
 sky130_fd_sc_hd__buf_6 _28772_ (.A(_19900_),
    .X(_06441_));
 sky130_fd_sc_hd__and4_2 _28773_ (.A(_19670_),
    .B(_05358_),
    .C(_06440_),
    .D(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__buf_8 _28774_ (.A(\pcpi_mul.rs1[15] ),
    .X(_06443_));
 sky130_fd_sc_hd__nand2_4 _28775_ (.A(_05290_),
    .B(_06443_),
    .Y(_06444_));
 sky130_vsdinv _28776_ (.A(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__o21ai_2 _28777_ (.A1(_06439_),
    .A2(_06442_),
    .B1(_06445_),
    .Y(_06446_));
 sky130_vsdinv _28778_ (.A(_05285_),
    .Y(_06447_));
 sky130_fd_sc_hd__buf_4 _28779_ (.A(_05642_),
    .X(_06448_));
 sky130_fd_sc_hd__nand2_1 _28780_ (.A(_05211_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__o21ai_2 _28781_ (.A1(_06447_),
    .A2(_05787_),
    .B1(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__nand3b_4 _28782_ (.A_N(_06449_),
    .B(_06258_),
    .C(_05977_),
    .Y(_06451_));
 sky130_fd_sc_hd__nand3_2 _28783_ (.A(_06450_),
    .B(_06451_),
    .C(_06444_),
    .Y(_06452_));
 sky130_fd_sc_hd__a21oi_2 _28784_ (.A1(_06273_),
    .A2(_06269_),
    .B1(_06266_),
    .Y(_06453_));
 sky130_fd_sc_hd__nand3_4 _28785_ (.A(_06446_),
    .B(_06452_),
    .C(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__nor2_2 _28786_ (.A(_06268_),
    .B(_06261_),
    .Y(_06455_));
 sky130_fd_sc_hd__nand3_2 _28787_ (.A(_06450_),
    .B(_06451_),
    .C(_06445_),
    .Y(_06456_));
 sky130_fd_sc_hd__o21ai_2 _28788_ (.A1(_06439_),
    .A2(_06442_),
    .B1(_06444_),
    .Y(_06457_));
 sky130_fd_sc_hd__o211ai_4 _28789_ (.A1(_06266_),
    .A2(_06455_),
    .B1(_06456_),
    .C1(_06457_),
    .Y(_06458_));
 sky130_vsdinv _28790_ (.A(_06287_),
    .Y(_06459_));
 sky130_fd_sc_hd__buf_4 _28791_ (.A(_06459_),
    .X(_06460_));
 sky130_fd_sc_hd__nor2_2 _28792_ (.A(_05132_),
    .B(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__buf_8 _28793_ (.A(_19890_),
    .X(_06462_));
 sky130_fd_sc_hd__a22oi_4 _28794_ (.A1(_05161_),
    .A2(_06462_),
    .B1(_05227_),
    .B2(_19888_),
    .Y(_06463_));
 sky130_fd_sc_hd__buf_6 _28795_ (.A(_19886_),
    .X(_06464_));
 sky130_fd_sc_hd__buf_6 _28796_ (.A(_06282_),
    .X(_06465_));
 sky130_fd_sc_hd__and4_2 _28797_ (.A(_05125_),
    .B(_19682_),
    .C(_06464_),
    .D(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__nor2_2 _28798_ (.A(_06463_),
    .B(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__nor2_2 _28799_ (.A(_06461_),
    .B(_06467_),
    .Y(_06468_));
 sky130_fd_sc_hd__and2_2 _28800_ (.A(_06467_),
    .B(_06461_),
    .X(_06469_));
 sky130_fd_sc_hd__o2bb2ai_4 _28801_ (.A1_N(_06454_),
    .A2_N(_06458_),
    .B1(_06468_),
    .B2(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__buf_6 _28802_ (.A(_06459_),
    .X(_06471_));
 sky130_fd_sc_hd__o21ai_1 _28803_ (.A1(_05491_),
    .A2(_06471_),
    .B1(_06467_),
    .Y(_06472_));
 sky130_fd_sc_hd__o21ai_1 _28804_ (.A1(_06463_),
    .A2(_06466_),
    .B1(_06461_),
    .Y(_06473_));
 sky130_fd_sc_hd__nand2_2 _28805_ (.A(_06472_),
    .B(_06473_),
    .Y(_06474_));
 sky130_fd_sc_hd__nand3_4 _28806_ (.A(_06474_),
    .B(_06458_),
    .C(_06454_),
    .Y(_06475_));
 sky130_fd_sc_hd__nand2_4 _28807_ (.A(_06303_),
    .B(_06279_),
    .Y(_06476_));
 sky130_fd_sc_hd__a21o_2 _28808_ (.A1(_06470_),
    .A2(_06475_),
    .B1(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__nand3_4 _28809_ (.A(_06476_),
    .B(_06470_),
    .C(_06475_),
    .Y(_06478_));
 sky130_fd_sc_hd__nor2_4 _28810_ (.A(_06290_),
    .B(_06291_),
    .Y(_06479_));
 sky130_vsdinv _28811_ (.A(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__nand3_4 _28812_ (.A(_06477_),
    .B(_06478_),
    .C(_06480_),
    .Y(_06481_));
 sky130_vsdinv _28813_ (.A(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__a21oi_2 _28814_ (.A1(_06477_),
    .A2(_06478_),
    .B1(_06480_),
    .Y(_06483_));
 sky130_vsdinv _28815_ (.A(_06232_),
    .Y(_06484_));
 sky130_fd_sc_hd__o21ai_4 _28816_ (.A1(_06078_),
    .A2(_06233_),
    .B1(_06227_),
    .Y(_06485_));
 sky130_vsdinv _28817_ (.A(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__a22oi_4 _28818_ (.A1(_05837_),
    .A2(_05666_),
    .B1(_19665_),
    .B2(_06106_),
    .Y(_06487_));
 sky130_fd_sc_hd__buf_4 _28819_ (.A(_05403_),
    .X(_06488_));
 sky130_fd_sc_hd__and4_4 _28820_ (.A(_19662_),
    .B(_06488_),
    .C(_19907_),
    .D(_05489_),
    .X(_06489_));
 sky130_fd_sc_hd__o22ai_4 _28821_ (.A1(_05261_),
    .A2(_05981_),
    .B1(_06487_),
    .B2(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__o21ai_2 _28822_ (.A1(_06333_),
    .A2(_06328_),
    .B1(_06337_),
    .Y(_06491_));
 sky130_fd_sc_hd__buf_4 _28823_ (.A(_05439_),
    .X(_06492_));
 sky130_fd_sc_hd__buf_8 _28824_ (.A(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__buf_6 _28825_ (.A(_05801_),
    .X(_06494_));
 sky130_fd_sc_hd__nand2_4 _28826_ (.A(_05699_),
    .B(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__a41oi_4 _28827_ (.A1(_06493_),
    .A2(_05405_),
    .A3(_05808_),
    .A4(_19911_),
    .B1(_06495_),
    .Y(_06496_));
 sky130_fd_sc_hd__a22o_1 _28828_ (.A1(_05587_),
    .A2(_05666_),
    .B1(_05589_),
    .B2(_06106_),
    .X(_06497_));
 sky130_fd_sc_hd__nand2_2 _28829_ (.A(_06496_),
    .B(_06497_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand3_4 _28830_ (.A(_06490_),
    .B(_06491_),
    .C(_06498_),
    .Y(_06499_));
 sky130_vsdinv _28831_ (.A(_06495_),
    .Y(_06500_));
 sky130_fd_sc_hd__o21ai_2 _28832_ (.A1(_06487_),
    .A2(_06489_),
    .B1(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__buf_6 _28833_ (.A(_19661_),
    .X(_06502_));
 sky130_fd_sc_hd__nand2_1 _28834_ (.A(_06502_),
    .B(_05770_),
    .Y(_06503_));
 sky130_fd_sc_hd__buf_6 _28835_ (.A(_06216_),
    .X(_06504_));
 sky130_fd_sc_hd__buf_8 _28836_ (.A(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__nand3b_4 _28837_ (.A_N(_06503_),
    .B(_06505_),
    .C(_19908_),
    .Y(_06506_));
 sky130_fd_sc_hd__nand3_4 _28838_ (.A(_06506_),
    .B(_06495_),
    .C(_06497_),
    .Y(_06507_));
 sky130_fd_sc_hd__o21ai_1 _28839_ (.A1(_06329_),
    .A2(_06331_),
    .B1(_06333_),
    .Y(_06508_));
 sky130_fd_sc_hd__nand2_1 _28840_ (.A(_06508_),
    .B(_06338_),
    .Y(_06509_));
 sky130_fd_sc_hd__nand3_4 _28841_ (.A(_06501_),
    .B(_06507_),
    .C(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__nor2_8 _28842_ (.A(_06222_),
    .B(_06219_),
    .Y(_06511_));
 sky130_fd_sc_hd__o2bb2ai_4 _28843_ (.A1_N(_06499_),
    .A2_N(_06510_),
    .B1(_06213_),
    .B2(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__nor2_4 _28844_ (.A(_06213_),
    .B(_06511_),
    .Y(_06513_));
 sky130_fd_sc_hd__nand3_4 _28845_ (.A(_06510_),
    .B(_06499_),
    .C(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__nand2_1 _28846_ (.A(_06360_),
    .B(_06340_),
    .Y(_06515_));
 sky130_fd_sc_hd__nand2_4 _28847_ (.A(_06515_),
    .B(_06357_),
    .Y(_06516_));
 sky130_fd_sc_hd__a21oi_4 _28848_ (.A1(_06512_),
    .A2(_06514_),
    .B1(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__and3_1 _28849_ (.A(_06490_),
    .B(_06491_),
    .C(_06498_),
    .X(_06518_));
 sky130_fd_sc_hd__nand2_1 _28850_ (.A(_06510_),
    .B(_06513_),
    .Y(_06519_));
 sky130_fd_sc_hd__o211a_2 _28851_ (.A1(_06518_),
    .A2(_06519_),
    .B1(_06512_),
    .C1(_06516_),
    .X(_06520_));
 sky130_fd_sc_hd__o22ai_4 _28852_ (.A1(_06484_),
    .A2(_06486_),
    .B1(_06517_),
    .B2(_06520_),
    .Y(_06521_));
 sky130_fd_sc_hd__nand2_4 _28853_ (.A(_06485_),
    .B(_06232_),
    .Y(_06522_));
 sky130_fd_sc_hd__a2bb2oi_2 _28854_ (.A1_N(_06213_),
    .A2_N(_06511_),
    .B1(_06499_),
    .B2(_06510_),
    .Y(_06523_));
 sky130_fd_sc_hd__nor2_1 _28855_ (.A(_06220_),
    .B(_06213_),
    .Y(_06524_));
 sky130_fd_sc_hd__o211a_1 _28856_ (.A1(_06219_),
    .A2(_06524_),
    .B1(_06499_),
    .C1(_06510_),
    .X(_06525_));
 sky130_fd_sc_hd__a21boi_4 _28857_ (.A1(_06360_),
    .A2(_06340_),
    .B1_N(_06357_),
    .Y(_06526_));
 sky130_fd_sc_hd__o21ai_4 _28858_ (.A1(_06523_),
    .A2(_06525_),
    .B1(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__nand3_4 _28859_ (.A(_06516_),
    .B(_06512_),
    .C(_06514_),
    .Y(_06528_));
 sky130_fd_sc_hd__nand3b_4 _28860_ (.A_N(_06522_),
    .B(_06527_),
    .C(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__o21ai_4 _28861_ (.A1(_06243_),
    .A2(_06237_),
    .B1(_06249_),
    .Y(_06530_));
 sky130_fd_sc_hd__a21oi_4 _28862_ (.A1(_06521_),
    .A2(_06529_),
    .B1(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__a21oi_1 _28863_ (.A1(_06246_),
    .A2(_06247_),
    .B1(_06243_),
    .Y(_06532_));
 sky130_fd_sc_hd__o211a_2 _28864_ (.A1(_06240_),
    .A2(_06532_),
    .B1(_06529_),
    .C1(_06521_),
    .X(_06533_));
 sky130_fd_sc_hd__o22ai_4 _28865_ (.A1(_06482_),
    .A2(_06483_),
    .B1(_06531_),
    .B2(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__and2_1 _28866_ (.A(_06249_),
    .B(_06243_),
    .X(_06535_));
 sky130_fd_sc_hd__a22oi_4 _28867_ (.A1(_06232_),
    .A2(_06485_),
    .B1(_06527_),
    .B2(_06528_),
    .Y(_06536_));
 sky130_fd_sc_hd__nor3_4 _28868_ (.A(_06522_),
    .B(_06517_),
    .C(_06520_),
    .Y(_06537_));
 sky130_fd_sc_hd__o22ai_4 _28869_ (.A1(_06237_),
    .A2(_06535_),
    .B1(_06536_),
    .B2(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__nand3_4 _28870_ (.A(_06521_),
    .B(_06530_),
    .C(_06529_),
    .Y(_06539_));
 sky130_fd_sc_hd__a21oi_4 _28871_ (.A1(_06470_),
    .A2(_06475_),
    .B1(_06476_),
    .Y(_06540_));
 sky130_fd_sc_hd__a32oi_4 _28872_ (.A1(_06270_),
    .A2(_06271_),
    .A3(_06274_),
    .B1(_06295_),
    .B2(_06296_),
    .Y(_06541_));
 sky130_fd_sc_hd__o211a_2 _28873_ (.A1(_06302_),
    .A2(_06541_),
    .B1(_06475_),
    .C1(_06470_),
    .X(_06542_));
 sky130_fd_sc_hd__o21ai_2 _28874_ (.A1(_06540_),
    .A2(_06542_),
    .B1(_06480_),
    .Y(_06543_));
 sky130_fd_sc_hd__nand3_2 _28875_ (.A(_06477_),
    .B(_06478_),
    .C(_06479_),
    .Y(_06544_));
 sky130_fd_sc_hd__nand2_4 _28876_ (.A(_06543_),
    .B(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__nand3_4 _28877_ (.A(_06538_),
    .B(_06539_),
    .C(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__nand2_1 _28878_ (.A(_06312_),
    .B(_06256_),
    .Y(_06547_));
 sky130_fd_sc_hd__nand2_4 _28879_ (.A(_06547_),
    .B(_06251_),
    .Y(_06548_));
 sky130_fd_sc_hd__a21oi_2 _28880_ (.A1(_06534_),
    .A2(_06546_),
    .B1(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__nand2_1 _28881_ (.A(_06538_),
    .B(_06545_),
    .Y(_06550_));
 sky130_fd_sc_hd__o211a_4 _28882_ (.A1(_06533_),
    .A2(_06550_),
    .B1(_06548_),
    .C1(_06534_),
    .X(_06551_));
 sky130_fd_sc_hd__o22ai_4 _28883_ (.A1(_06437_),
    .A2(_06438_),
    .B1(_06549_),
    .B2(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__o21ai_2 _28884_ (.A1(_06540_),
    .A2(_06542_),
    .B1(_06479_),
    .Y(_06553_));
 sky130_fd_sc_hd__a22oi_4 _28885_ (.A1(_06481_),
    .A2(_06553_),
    .B1(_06538_),
    .B2(_06539_),
    .Y(_06554_));
 sky130_fd_sc_hd__nand2_2 _28886_ (.A(_06521_),
    .B(_06530_),
    .Y(_06555_));
 sky130_fd_sc_hd__o211a_1 _28887_ (.A1(_06537_),
    .A2(_06555_),
    .B1(_06545_),
    .C1(_06538_),
    .X(_06556_));
 sky130_fd_sc_hd__o21bai_4 _28888_ (.A1(_06554_),
    .A2(_06556_),
    .B1_N(_06548_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand3_4 _28889_ (.A(_06534_),
    .B(_06548_),
    .C(_06546_),
    .Y(_06558_));
 sky130_fd_sc_hd__nor2_4 _28890_ (.A(_06438_),
    .B(_06437_),
    .Y(_06559_));
 sky130_fd_sc_hd__nand3_4 _28891_ (.A(_06557_),
    .B(_06558_),
    .C(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__a22oi_4 _28892_ (.A1(_06369_),
    .A2(_06325_),
    .B1(_06552_),
    .B2(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__nand2_2 _28893_ (.A(_06557_),
    .B(_06559_),
    .Y(_06562_));
 sky130_fd_sc_hd__o211a_1 _28894_ (.A1(_06551_),
    .A2(_06562_),
    .B1(_06372_),
    .C1(_06552_),
    .X(_06563_));
 sky130_fd_sc_hd__o22ai_4 _28895_ (.A1(_06396_),
    .A2(_06397_),
    .B1(_06561_),
    .B2(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__a21o_1 _28896_ (.A1(_06552_),
    .A2(_06560_),
    .B1(_06372_),
    .X(_06565_));
 sky130_fd_sc_hd__nand3_4 _28897_ (.A(_06552_),
    .B(_06372_),
    .C(_06560_),
    .Y(_06566_));
 sky130_fd_sc_hd__nor2_8 _28898_ (.A(_06397_),
    .B(_06396_),
    .Y(_06567_));
 sky130_fd_sc_hd__nand3_2 _28899_ (.A(_06565_),
    .B(_06566_),
    .C(_06567_),
    .Y(_06568_));
 sky130_fd_sc_hd__a22oi_4 _28900_ (.A1(_06366_),
    .A2(_06370_),
    .B1(_06373_),
    .B2(_06212_),
    .Y(_06569_));
 sky130_fd_sc_hd__nand3_4 _28901_ (.A(_06564_),
    .B(_06568_),
    .C(_06569_),
    .Y(_06570_));
 sky130_fd_sc_hd__o211a_1 _28902_ (.A1(_06396_),
    .A2(_06397_),
    .B1(_06566_),
    .C1(_06565_),
    .X(_06571_));
 sky130_fd_sc_hd__nand2_1 _28903_ (.A(_06373_),
    .B(_06212_),
    .Y(_06572_));
 sky130_fd_sc_hd__nand2_1 _28904_ (.A(_06572_),
    .B(_06371_),
    .Y(_06573_));
 sky130_fd_sc_hd__o21ai_1 _28905_ (.A1(_06561_),
    .A2(_06563_),
    .B1(_06567_),
    .Y(_06574_));
 sky130_fd_sc_hd__nand2_1 _28906_ (.A(_06573_),
    .B(_06574_),
    .Y(_06575_));
 sky130_fd_sc_hd__or2_1 _28907_ (.A(_06571_),
    .B(_06575_),
    .X(_06576_));
 sky130_fd_sc_hd__a21o_1 _28908_ (.A1(_06576_),
    .A2(_06570_),
    .B1(_06210_),
    .X(_06577_));
 sky130_fd_sc_hd__a21boi_4 _28909_ (.A1(_06210_),
    .A2(_06570_),
    .B1_N(_06577_),
    .Y(_06578_));
 sky130_fd_sc_hd__or2_1 _28910_ (.A(_06393_),
    .B(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__nand2_2 _28911_ (.A(_06385_),
    .B(_06379_),
    .Y(_06580_));
 sky130_fd_sc_hd__nand2_1 _28912_ (.A(_06392_),
    .B(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__nand2_1 _28913_ (.A(_06578_),
    .B(_06393_),
    .Y(_06582_));
 sky130_fd_sc_hd__nand3_4 _28914_ (.A(_06392_),
    .B(_06580_),
    .C(_06582_),
    .Y(_06583_));
 sky130_fd_sc_hd__and2_4 _28915_ (.A(_06583_),
    .B(_06579_),
    .X(_06584_));
 sky130_vsdinv _28916_ (.A(_06584_),
    .Y(_06585_));
 sky130_fd_sc_hd__o21a_1 _28917_ (.A1(_06579_),
    .A2(_06581_),
    .B1(_06585_),
    .X(_02634_));
 sky130_fd_sc_hd__a21oi_4 _28918_ (.A1(_06477_),
    .A2(_06480_),
    .B1(_06542_),
    .Y(_06586_));
 sky130_fd_sc_hd__nor2_4 _28919_ (.A(_06586_),
    .B(_06558_),
    .Y(_06587_));
 sky130_fd_sc_hd__and2_1 _28920_ (.A(_06558_),
    .B(_06586_),
    .X(_06588_));
 sky130_fd_sc_hd__nor2_4 _28921_ (.A(_06587_),
    .B(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__nand2_1 _28922_ (.A(_19637_),
    .B(_19934_),
    .Y(_06590_));
 sky130_fd_sc_hd__nand2_1 _28923_ (.A(net458),
    .B(_19931_),
    .Y(_06591_));
 sky130_fd_sc_hd__nand2_1 _28924_ (.A(_06590_),
    .B(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__or2_4 _28925_ (.A(_06590_),
    .B(_06591_),
    .X(_06593_));
 sky130_fd_sc_hd__nand2_1 _28926_ (.A(_06022_),
    .B(_05268_),
    .Y(_06594_));
 sky130_fd_sc_hd__nand2_1 _28927_ (.A(_05736_),
    .B(_05656_),
    .Y(_06595_));
 sky130_fd_sc_hd__nor2_2 _28928_ (.A(_06594_),
    .B(_06595_),
    .Y(_06596_));
 sky130_fd_sc_hd__nand2_2 _28929_ (.A(_19659_),
    .B(_05489_),
    .Y(_06597_));
 sky130_fd_sc_hd__nand2_1 _28930_ (.A(_06594_),
    .B(_06595_),
    .Y(_06598_));
 sky130_fd_sc_hd__nand3b_1 _28931_ (.A_N(_06596_),
    .B(_06597_),
    .C(_06598_),
    .Y(_06599_));
 sky130_fd_sc_hd__a22oi_4 _28932_ (.A1(net477),
    .A2(_05493_),
    .B1(_06399_),
    .B2(_19914_),
    .Y(_06600_));
 sky130_vsdinv _28933_ (.A(_06597_),
    .Y(_06601_));
 sky130_fd_sc_hd__o21ai_1 _28934_ (.A1(_06600_),
    .A2(_06596_),
    .B1(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__nand2_2 _28935_ (.A(_06599_),
    .B(_06602_),
    .Y(_06603_));
 sky130_vsdinv _28936_ (.A(_06603_),
    .Y(_06604_));
 sky130_fd_sc_hd__buf_4 _28937_ (.A(\pcpi_mul.rs2[14] ),
    .X(_06605_));
 sky130_fd_sc_hd__buf_6 _28938_ (.A(_06605_),
    .X(_06606_));
 sky130_fd_sc_hd__a22oi_4 _28939_ (.A1(_06606_),
    .A2(_05128_),
    .B1(_06169_),
    .B2(_06015_),
    .Y(_06607_));
 sky130_fd_sc_hd__buf_8 _28940_ (.A(_06413_),
    .X(_06608_));
 sky130_fd_sc_hd__nand2_2 _28941_ (.A(_06608_),
    .B(_05127_),
    .Y(_06609_));
 sky130_fd_sc_hd__buf_6 _28942_ (.A(_06167_),
    .X(_06610_));
 sky130_fd_sc_hd__nand2_2 _28943_ (.A(_06610_),
    .B(_05359_),
    .Y(_06611_));
 sky130_fd_sc_hd__nor2_4 _28944_ (.A(_06609_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__nand2_2 _28945_ (.A(_06419_),
    .B(_19920_),
    .Y(_06613_));
 sky130_fd_sc_hd__o21a_1 _28946_ (.A1(_06607_),
    .A2(_06612_),
    .B1(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__o21ai_2 _28947_ (.A1(_06415_),
    .A2(_06417_),
    .B1(_06420_),
    .Y(_06615_));
 sky130_fd_sc_hd__o311ai_4 _28948_ (.A1(_06613_),
    .A2(_06607_),
    .A3(_06612_),
    .B1(_06425_),
    .C1(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__o21bai_2 _28949_ (.A1(_06607_),
    .A2(_06612_),
    .B1_N(_06613_),
    .Y(_06617_));
 sky130_fd_sc_hd__clkbuf_8 _28950_ (.A(_19647_),
    .X(_06618_));
 sky130_fd_sc_hd__nand3b_1 _28951_ (.A_N(_06609_),
    .B(_06618_),
    .C(_19925_),
    .Y(_06619_));
 sky130_fd_sc_hd__nand2_1 _28952_ (.A(_06609_),
    .B(_06611_),
    .Y(_06620_));
 sky130_fd_sc_hd__nand3_2 _28953_ (.A(_06619_),
    .B(_06613_),
    .C(_06620_),
    .Y(_06621_));
 sky130_fd_sc_hd__nand2_1 _28954_ (.A(_06615_),
    .B(_06425_),
    .Y(_06622_));
 sky130_fd_sc_hd__nand3_4 _28955_ (.A(_06617_),
    .B(_06621_),
    .C(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__o21ai_2 _28956_ (.A1(_06614_),
    .A2(_06616_),
    .B1(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__or2_2 _28957_ (.A(_06604_),
    .B(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__nand2_2 _28958_ (.A(_06624_),
    .B(_06604_),
    .Y(_06626_));
 sky130_fd_sc_hd__a22o_2 _28959_ (.A1(_06592_),
    .A2(_06593_),
    .B1(_06625_),
    .B2(_06626_),
    .X(_06627_));
 sky130_fd_sc_hd__nand2_1 _28960_ (.A(_06593_),
    .B(_06592_),
    .Y(_06628_));
 sky130_fd_sc_hd__nand3b_4 _28961_ (.A_N(_06628_),
    .B(_06625_),
    .C(_06626_),
    .Y(_06629_));
 sky130_fd_sc_hd__nand2_4 _28962_ (.A(_06627_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__nor2_4 _28963_ (.A(_06436_),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__and2_1 _28964_ (.A(_06630_),
    .B(_06436_),
    .X(_06632_));
 sky130_fd_sc_hd__nand2_1 _28965_ (.A(_06475_),
    .B(_06458_),
    .Y(_06633_));
 sky130_fd_sc_hd__buf_4 _28966_ (.A(\pcpi_mul.rs1[15] ),
    .X(_06634_));
 sky130_fd_sc_hd__buf_4 _28967_ (.A(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__clkbuf_4 _28968_ (.A(_05116_),
    .X(_06636_));
 sky130_fd_sc_hd__nand2_2 _28969_ (.A(_06636_),
    .B(_19888_),
    .Y(_06637_));
 sky130_fd_sc_hd__a21o_2 _28970_ (.A1(_05235_),
    .A2(_06635_),
    .B1(_06637_),
    .X(_06638_));
 sky130_fd_sc_hd__buf_4 _28971_ (.A(_05266_),
    .X(_06639_));
 sky130_fd_sc_hd__buf_6 _28972_ (.A(_06267_),
    .X(_06640_));
 sky130_fd_sc_hd__buf_4 _28973_ (.A(_19883_),
    .X(_06641_));
 sky130_fd_sc_hd__nand2_2 _28974_ (.A(_05163_),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__a21o_2 _28975_ (.A1(_06639_),
    .A2(_06640_),
    .B1(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__nand2_2 _28976_ (.A(_05157_),
    .B(_19892_),
    .Y(_06644_));
 sky130_fd_sc_hd__a21oi_4 _28977_ (.A1(_06638_),
    .A2(_06643_),
    .B1(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__nand3_2 _28978_ (.A(_06638_),
    .B(_06643_),
    .C(_06644_),
    .Y(_06646_));
 sky130_fd_sc_hd__and2b_1 _28979_ (.A_N(_06645_),
    .B(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__buf_6 _28980_ (.A(_06117_),
    .X(_06648_));
 sky130_fd_sc_hd__buf_6 _28981_ (.A(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__clkbuf_8 _28982_ (.A(_06115_),
    .X(_06650_));
 sky130_fd_sc_hd__a22oi_4 _28983_ (.A1(_05778_),
    .A2(_06649_),
    .B1(_06258_),
    .B2(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__buf_6 _28984_ (.A(_06287_),
    .X(_06652_));
 sky130_fd_sc_hd__and4_2 _28985_ (.A(_05772_),
    .B(_05282_),
    .C(_06652_),
    .D(_19898_),
    .X(_06653_));
 sky130_fd_sc_hd__buf_8 _28986_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06654_));
 sky130_fd_sc_hd__nand2_4 _28987_ (.A(net495),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__o21ai_4 _28988_ (.A1(_06651_),
    .A2(_06653_),
    .B1(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__buf_4 _28989_ (.A(_06117_),
    .X(_06657_));
 sky130_fd_sc_hd__nand2_1 _28990_ (.A(_19670_),
    .B(_06657_),
    .Y(_06658_));
 sky130_fd_sc_hd__buf_6 _28991_ (.A(_05285_),
    .X(_06659_));
 sky130_fd_sc_hd__nand3b_4 _28992_ (.A_N(_06658_),
    .B(_06659_),
    .C(_06289_),
    .Y(_06660_));
 sky130_vsdinv _28993_ (.A(_06655_),
    .Y(_06661_));
 sky130_fd_sc_hd__a22o_2 _28994_ (.A1(_05295_),
    .A2(_06649_),
    .B1(_19673_),
    .B2(_06650_),
    .X(_06662_));
 sky130_fd_sc_hd__nand3_4 _28995_ (.A(_06660_),
    .B(_06661_),
    .C(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__o21ai_4 _28996_ (.A1(_06444_),
    .A2(_06439_),
    .B1(_06451_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand3_4 _28997_ (.A(_06656_),
    .B(_06663_),
    .C(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__o21ai_2 _28998_ (.A1(_06651_),
    .A2(_06653_),
    .B1(_06661_),
    .Y(_06666_));
 sky130_fd_sc_hd__nand3_2 _28999_ (.A(_06660_),
    .B(_06655_),
    .C(_06662_),
    .Y(_06667_));
 sky130_fd_sc_hd__nand3b_4 _29000_ (.A_N(_06664_),
    .B(_06666_),
    .C(_06667_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand3_2 _29001_ (.A(_06647_),
    .B(_06665_),
    .C(_06668_),
    .Y(_06669_));
 sky130_fd_sc_hd__nand2_1 _29002_ (.A(_06668_),
    .B(_06665_),
    .Y(_06670_));
 sky130_fd_sc_hd__a21o_1 _29003_ (.A1(_06638_),
    .A2(_06643_),
    .B1(_06644_),
    .X(_06671_));
 sky130_fd_sc_hd__nand2_2 _29004_ (.A(_06671_),
    .B(_06646_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand2_1 _29005_ (.A(_06670_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nand3_4 _29006_ (.A(_06633_),
    .B(_06669_),
    .C(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__nand2_1 _29007_ (.A(_06670_),
    .B(_06647_),
    .Y(_06675_));
 sky130_fd_sc_hd__a21boi_2 _29008_ (.A1(_06474_),
    .A2(_06454_),
    .B1_N(_06458_),
    .Y(_06676_));
 sky130_fd_sc_hd__nand3_2 _29009_ (.A(_06672_),
    .B(_06668_),
    .C(_06665_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand3_4 _29010_ (.A(_06675_),
    .B(_06676_),
    .C(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__nor2_4 _29011_ (.A(_06466_),
    .B(_06469_),
    .Y(_06679_));
 sky130_vsdinv _29012_ (.A(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__and3_4 _29013_ (.A(_06674_),
    .B(_06678_),
    .C(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__a21oi_4 _29014_ (.A1(_06674_),
    .A2(_06678_),
    .B1(_06680_),
    .Y(_06682_));
 sky130_fd_sc_hd__nand2_1 _29015_ (.A(_06528_),
    .B(_06522_),
    .Y(_06683_));
 sky130_vsdinv _29016_ (.A(_06510_),
    .Y(_06684_));
 sky130_fd_sc_hd__nor2_2 _29017_ (.A(_06513_),
    .B(_06518_),
    .Y(_06685_));
 sky130_fd_sc_hd__buf_6 _29018_ (.A(_05464_),
    .X(_06686_));
 sky130_fd_sc_hd__a22oi_4 _29019_ (.A1(_06076_),
    .A2(_06686_),
    .B1(_06077_),
    .B2(_05797_),
    .Y(_06687_));
 sky130_fd_sc_hd__nand3_4 _29020_ (.A(_05451_),
    .B(_06217_),
    .C(_05958_),
    .Y(_06688_));
 sky130_fd_sc_hd__nor2_8 _29021_ (.A(net447),
    .B(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__nand2_1 _29022_ (.A(_05835_),
    .B(_06441_),
    .Y(_06690_));
 sky130_vsdinv _29023_ (.A(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__o21bai_2 _29024_ (.A1(_06687_),
    .A2(_06689_),
    .B1_N(_06691_),
    .Y(_06692_));
 sky130_fd_sc_hd__o21ai_2 _29025_ (.A1(_06405_),
    .A2(_06400_),
    .B1(_06407_),
    .Y(_06693_));
 sky130_fd_sc_hd__a22o_2 _29026_ (.A1(_05587_),
    .A2(_06686_),
    .B1(_05589_),
    .B2(_05797_),
    .X(_06694_));
 sky130_fd_sc_hd__o211ai_4 _29027_ (.A1(_05981_),
    .A2(_06688_),
    .B1(_06691_),
    .C1(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__nand3_4 _29028_ (.A(_06692_),
    .B(_06693_),
    .C(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__o21ai_2 _29029_ (.A1(_06687_),
    .A2(_06689_),
    .B1(_06691_),
    .Y(_06697_));
 sky130_fd_sc_hd__o21ai_1 _29030_ (.A1(_06402_),
    .A2(_06403_),
    .B1(_06405_),
    .Y(_06698_));
 sky130_fd_sc_hd__nand2_1 _29031_ (.A(_06698_),
    .B(_06408_),
    .Y(_06699_));
 sky130_fd_sc_hd__o211ai_2 _29032_ (.A1(_05981_),
    .A2(_06688_),
    .B1(_06690_),
    .C1(_06694_),
    .Y(_06700_));
 sky130_fd_sc_hd__nand3_4 _29033_ (.A(_06697_),
    .B(_06699_),
    .C(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__nor2_4 _29034_ (.A(_06500_),
    .B(_06489_),
    .Y(_06702_));
 sky130_fd_sc_hd__o2bb2ai_4 _29035_ (.A1_N(_06696_),
    .A2_N(_06701_),
    .B1(_06487_),
    .B2(_06702_),
    .Y(_06703_));
 sky130_fd_sc_hd__nor2_4 _29036_ (.A(_06487_),
    .B(_06702_),
    .Y(_06704_));
 sky130_fd_sc_hd__nand3_4 _29037_ (.A(_06701_),
    .B(_06696_),
    .C(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__nand2_1 _29038_ (.A(_06430_),
    .B(_06410_),
    .Y(_06706_));
 sky130_fd_sc_hd__nand2_4 _29039_ (.A(_06706_),
    .B(_06429_),
    .Y(_06707_));
 sky130_fd_sc_hd__a21oi_4 _29040_ (.A1(_06703_),
    .A2(_06705_),
    .B1(_06707_),
    .Y(_06708_));
 sky130_fd_sc_hd__and3_1 _29041_ (.A(_06692_),
    .B(_06693_),
    .C(_06695_),
    .X(_06709_));
 sky130_fd_sc_hd__nand2_1 _29042_ (.A(_06701_),
    .B(_06704_),
    .Y(_06710_));
 sky130_fd_sc_hd__o211a_2 _29043_ (.A1(_06709_),
    .A2(_06710_),
    .B1(_06703_),
    .C1(_06707_),
    .X(_06711_));
 sky130_fd_sc_hd__o22ai_4 _29044_ (.A1(_06684_),
    .A2(_06685_),
    .B1(_06708_),
    .B2(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__nand2_1 _29045_ (.A(_06703_),
    .B(_06705_),
    .Y(_06713_));
 sky130_fd_sc_hd__and2_1 _29046_ (.A(_06706_),
    .B(_06429_),
    .X(_06714_));
 sky130_fd_sc_hd__nand2_1 _29047_ (.A(_06713_),
    .B(_06714_),
    .Y(_06715_));
 sky130_fd_sc_hd__nand3_4 _29048_ (.A(_06707_),
    .B(_06703_),
    .C(_06705_),
    .Y(_06716_));
 sky130_fd_sc_hd__nand2_2 _29049_ (.A(_06519_),
    .B(_06499_),
    .Y(_06717_));
 sky130_fd_sc_hd__nand3_4 _29050_ (.A(_06715_),
    .B(_06716_),
    .C(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__a22oi_4 _29051_ (.A1(_06527_),
    .A2(_06683_),
    .B1(_06712_),
    .B2(_06718_),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_1 _29052_ (.A(_06512_),
    .B(_06514_),
    .Y(_06720_));
 sky130_fd_sc_hd__a21oi_1 _29053_ (.A1(_06720_),
    .A2(_06526_),
    .B1(_06522_),
    .Y(_06721_));
 sky130_fd_sc_hd__o211a_4 _29054_ (.A1(_06520_),
    .A2(_06721_),
    .B1(_06718_),
    .C1(_06712_),
    .X(_06722_));
 sky130_fd_sc_hd__o22ai_4 _29055_ (.A1(_06681_),
    .A2(_06682_),
    .B1(_06719_),
    .B2(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__nand2_1 _29056_ (.A(_06553_),
    .B(_06481_),
    .Y(_06724_));
 sky130_fd_sc_hd__o22ai_4 _29057_ (.A1(_06537_),
    .A2(_06555_),
    .B1(_06724_),
    .B2(_06531_),
    .Y(_06725_));
 sky130_fd_sc_hd__o21ai_2 _29058_ (.A1(_06522_),
    .A2(_06517_),
    .B1(_06528_),
    .Y(_06726_));
 sky130_fd_sc_hd__a21o_1 _29059_ (.A1(_06712_),
    .A2(_06718_),
    .B1(_06726_),
    .X(_06727_));
 sky130_fd_sc_hd__nand3_4 _29060_ (.A(_06712_),
    .B(_06726_),
    .C(_06718_),
    .Y(_06728_));
 sky130_fd_sc_hd__nor2_8 _29061_ (.A(_06682_),
    .B(_06681_),
    .Y(_06729_));
 sky130_fd_sc_hd__nand3_4 _29062_ (.A(_06727_),
    .B(_06728_),
    .C(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__nand3_4 _29063_ (.A(_06723_),
    .B(_06725_),
    .C(_06730_),
    .Y(_06731_));
 sky130_fd_sc_hd__clkbuf_4 _29064_ (.A(_06731_),
    .X(_06732_));
 sky130_fd_sc_hd__o21ai_2 _29065_ (.A1(_06719_),
    .A2(_06722_),
    .B1(_06729_),
    .Y(_06733_));
 sky130_fd_sc_hd__a21oi_4 _29066_ (.A1(_06538_),
    .A2(_06545_),
    .B1(_06533_),
    .Y(_06734_));
 sky130_fd_sc_hd__a21o_1 _29067_ (.A1(_06674_),
    .A2(_06678_),
    .B1(_06680_),
    .X(_06735_));
 sky130_fd_sc_hd__nand3_1 _29068_ (.A(_06674_),
    .B(_06678_),
    .C(_06680_),
    .Y(_06736_));
 sky130_fd_sc_hd__nand2_1 _29069_ (.A(_06735_),
    .B(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__nand3_2 _29070_ (.A(_06727_),
    .B(_06728_),
    .C(_06737_),
    .Y(_06738_));
 sky130_fd_sc_hd__nand3_4 _29071_ (.A(_06733_),
    .B(_06734_),
    .C(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__a2bb2oi_2 _29072_ (.A1_N(_06631_),
    .A2_N(_06632_),
    .B1(_06732_),
    .B2(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__and2_2 _29073_ (.A(_06630_),
    .B(_06437_),
    .X(_06741_));
 sky130_fd_sc_hd__nor2_4 _29074_ (.A(_06437_),
    .B(_06630_),
    .Y(_06742_));
 sky130_fd_sc_hd__o211a_1 _29075_ (.A1(_06741_),
    .A2(_06742_),
    .B1(_06731_),
    .C1(_06739_),
    .X(_06743_));
 sky130_fd_sc_hd__o22ai_4 _29076_ (.A1(_06551_),
    .A2(_06562_),
    .B1(_06740_),
    .B2(_06743_),
    .Y(_06744_));
 sky130_vsdinv _29077_ (.A(_06548_),
    .Y(_06745_));
 sky130_fd_sc_hd__nand2_2 _29078_ (.A(_06534_),
    .B(_06546_),
    .Y(_06746_));
 sky130_fd_sc_hd__o211ai_4 _29079_ (.A1(_06741_),
    .A2(_06742_),
    .B1(_06731_),
    .C1(_06739_),
    .Y(_06747_));
 sky130_fd_sc_hd__a21boi_2 _29080_ (.A1(_06745_),
    .A2(_06746_),
    .B1_N(_06559_),
    .Y(_06748_));
 sky130_fd_sc_hd__o2bb2ai_1 _29081_ (.A1_N(_06732_),
    .A2_N(_06739_),
    .B1(_06631_),
    .B2(_06632_),
    .Y(_06749_));
 sky130_fd_sc_hd__o2111ai_4 _29082_ (.A1(_06745_),
    .A2(_06746_),
    .B1(_06747_),
    .C1(_06748_),
    .D1(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__nand3b_2 _29083_ (.A_N(_06589_),
    .B(_06744_),
    .C(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__nor2_1 _29084_ (.A(_06586_),
    .B(_06551_),
    .Y(_06752_));
 sky130_fd_sc_hd__and2_1 _29085_ (.A(_06551_),
    .B(_06586_),
    .X(_06753_));
 sky130_fd_sc_hd__o2bb2ai_1 _29086_ (.A1_N(_06750_),
    .A2_N(_06744_),
    .B1(_06752_),
    .B2(_06753_),
    .Y(_06754_));
 sky130_fd_sc_hd__o2111ai_4 _29087_ (.A1(_06561_),
    .A2(_06567_),
    .B1(_06566_),
    .C1(_06751_),
    .D1(_06754_),
    .Y(_06755_));
 sky130_vsdinv _29088_ (.A(_06560_),
    .Y(_06756_));
 sky130_fd_sc_hd__nand2_1 _29089_ (.A(_06552_),
    .B(_06372_),
    .Y(_06757_));
 sky130_fd_sc_hd__o22ai_4 _29090_ (.A1(_06756_),
    .A2(_06757_),
    .B1(_06567_),
    .B2(_06561_),
    .Y(_06758_));
 sky130_fd_sc_hd__o2bb2ai_1 _29091_ (.A1_N(_06750_),
    .A2_N(_06744_),
    .B1(_06587_),
    .B2(_06588_),
    .Y(_06759_));
 sky130_fd_sc_hd__nand3_2 _29092_ (.A(_06744_),
    .B(_06750_),
    .C(_06589_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand3_4 _29093_ (.A(_06758_),
    .B(_06759_),
    .C(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nor2_4 _29094_ (.A(_06394_),
    .B(_06325_),
    .Y(_06762_));
 sky130_fd_sc_hd__a21oi_1 _29095_ (.A1(_06755_),
    .A2(_06761_),
    .B1(_06762_),
    .Y(_06763_));
 sky130_fd_sc_hd__and3_1 _29096_ (.A(_06755_),
    .B(_06761_),
    .C(_06762_),
    .X(_06764_));
 sky130_fd_sc_hd__o2bb2ai_2 _29097_ (.A1_N(_06210_),
    .A2_N(_06570_),
    .B1(_06571_),
    .B2(_06575_),
    .Y(_06765_));
 sky130_fd_sc_hd__o21bai_2 _29098_ (.A1(_06763_),
    .A2(_06764_),
    .B1_N(_06765_),
    .Y(_06766_));
 sky130_fd_sc_hd__a21o_1 _29099_ (.A1(_06755_),
    .A2(_06761_),
    .B1(_06762_),
    .X(_06767_));
 sky130_fd_sc_hd__nand3_4 _29100_ (.A(_06755_),
    .B(_06761_),
    .C(_06762_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand3_4 _29101_ (.A(_06767_),
    .B(_06765_),
    .C(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__nand2_2 _29102_ (.A(_06766_),
    .B(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__and2_1 _29103_ (.A(_06585_),
    .B(_06770_),
    .X(_06771_));
 sky130_fd_sc_hd__a21oi_4 _29104_ (.A1(_06584_),
    .A2(_06766_),
    .B1(_06771_),
    .Y(_02635_));
 sky130_vsdinv _29105_ (.A(_06678_),
    .Y(_06772_));
 sky130_fd_sc_hd__a21oi_4 _29106_ (.A1(_06679_),
    .A2(_06674_),
    .B1(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__and2_2 _29107_ (.A(_06731_),
    .B(_06773_),
    .X(_06774_));
 sky130_fd_sc_hd__nor2_4 _29108_ (.A(_06773_),
    .B(_06732_),
    .Y(_06775_));
 sky130_fd_sc_hd__nand2_2 _29109_ (.A(_06739_),
    .B(_06732_),
    .Y(_06776_));
 sky130_fd_sc_hd__nor2_4 _29110_ (.A(_06742_),
    .B(_06741_),
    .Y(_06777_));
 sky130_fd_sc_hd__nor2_4 _29111_ (.A(_06637_),
    .B(_06642_),
    .Y(_06778_));
 sky130_fd_sc_hd__buf_4 _29112_ (.A(\pcpi_mul.rs1[13] ),
    .X(_06779_));
 sky130_fd_sc_hd__clkbuf_8 _29113_ (.A(_06779_),
    .X(_06780_));
 sky130_fd_sc_hd__a22oi_4 _29114_ (.A1(_05212_),
    .A2(_06116_),
    .B1(_06659_),
    .B2(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__and4_2 _29115_ (.A(_05212_),
    .B(_06258_),
    .C(_19891_),
    .D(_06116_),
    .X(_06782_));
 sky130_fd_sc_hd__clkbuf_8 _29116_ (.A(\pcpi_mul.rs1[17] ),
    .X(_06783_));
 sky130_fd_sc_hd__nand2_4 _29117_ (.A(_05290_),
    .B(_06783_),
    .Y(_06784_));
 sky130_vsdinv _29118_ (.A(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__o21ai_2 _29119_ (.A1(_06781_),
    .A2(_06782_),
    .B1(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__a21oi_2 _29120_ (.A1(_06662_),
    .A2(_06661_),
    .B1(_06653_),
    .Y(_06787_));
 sky130_fd_sc_hd__buf_8 _29121_ (.A(_19893_),
    .X(_06788_));
 sky130_fd_sc_hd__nand2_1 _29122_ (.A(_05197_),
    .B(_06788_),
    .Y(_06789_));
 sky130_fd_sc_hd__nand3b_4 _29123_ (.A_N(_06789_),
    .B(_05792_),
    .C(_06284_),
    .Y(_06790_));
 sky130_fd_sc_hd__a22o_1 _29124_ (.A1(_05212_),
    .A2(_06289_),
    .B1(_06659_),
    .B2(_06286_),
    .X(_06791_));
 sky130_fd_sc_hd__nand3_2 _29125_ (.A(_06790_),
    .B(_06791_),
    .C(_06784_),
    .Y(_06792_));
 sky130_fd_sc_hd__nand3_4 _29126_ (.A(_06786_),
    .B(_06787_),
    .C(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__o21ai_2 _29127_ (.A1(_06781_),
    .A2(_06782_),
    .B1(_06784_),
    .Y(_06794_));
 sky130_fd_sc_hd__nand3_2 _29128_ (.A(_06790_),
    .B(_06791_),
    .C(_06785_),
    .Y(_06795_));
 sky130_fd_sc_hd__o21ai_2 _29129_ (.A1(_06655_),
    .A2(_06651_),
    .B1(_06660_),
    .Y(_06796_));
 sky130_fd_sc_hd__nand3_4 _29130_ (.A(_06794_),
    .B(_06795_),
    .C(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__clkbuf_4 _29131_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06798_));
 sky130_fd_sc_hd__buf_6 _29132_ (.A(_06798_),
    .X(_06799_));
 sky130_fd_sc_hd__nand2_2 _29133_ (.A(_05227_),
    .B(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__nand3_4 _29134_ (.A(_06800_),
    .B(_06639_),
    .C(_06635_),
    .Y(_06801_));
 sky130_fd_sc_hd__nand2_2 _29135_ (.A(_19679_),
    .B(_06641_),
    .Y(_06802_));
 sky130_fd_sc_hd__clkbuf_8 _29136_ (.A(\pcpi_mul.rs1[16] ),
    .X(_06803_));
 sky130_fd_sc_hd__clkbuf_8 _29137_ (.A(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__nand3_4 _29138_ (.A(_06802_),
    .B(_05235_),
    .C(_06804_),
    .Y(_06805_));
 sky130_fd_sc_hd__nand2_1 _29139_ (.A(_05807_),
    .B(net435),
    .Y(_06806_));
 sky130_fd_sc_hd__a21oi_4 _29140_ (.A1(_06801_),
    .A2(_06805_),
    .B1(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__clkbuf_4 _29141_ (.A(\pcpi_mul.rs1[14] ),
    .X(_06808_));
 sky130_vsdinv _29142_ (.A(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__buf_6 _29143_ (.A(_06809_),
    .X(_06810_));
 sky130_fd_sc_hd__o211a_2 _29144_ (.A1(_05491_),
    .A2(_06810_),
    .B1(_06801_),
    .C1(_06805_),
    .X(_06811_));
 sky130_fd_sc_hd__nor2_8 _29145_ (.A(_06807_),
    .B(_06811_),
    .Y(_06812_));
 sky130_fd_sc_hd__a21oi_4 _29146_ (.A1(_06793_),
    .A2(_06797_),
    .B1(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__a21oi_4 _29147_ (.A1(_06656_),
    .A2(_06663_),
    .B1(_06664_),
    .Y(_06814_));
 sky130_fd_sc_hd__o21ai_2 _29148_ (.A1(_06814_),
    .A2(_06672_),
    .B1(_06665_),
    .Y(_06815_));
 sky130_fd_sc_hd__nand3_2 _29149_ (.A(_06812_),
    .B(_06793_),
    .C(_06797_),
    .Y(_06816_));
 sky130_fd_sc_hd__nand3b_4 _29150_ (.A_N(_06813_),
    .B(_06815_),
    .C(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__and3_1 _29151_ (.A(_06812_),
    .B(_06793_),
    .C(_06797_),
    .X(_06818_));
 sky130_fd_sc_hd__o21a_1 _29152_ (.A1(_06814_),
    .A2(_06672_),
    .B1(_06665_),
    .X(_06819_));
 sky130_fd_sc_hd__o21ai_4 _29153_ (.A1(_06813_),
    .A2(_06818_),
    .B1(_06819_),
    .Y(_06820_));
 sky130_fd_sc_hd__o211a_2 _29154_ (.A1(_06778_),
    .A2(_06645_),
    .B1(_06817_),
    .C1(_06820_),
    .X(_06821_));
 sky130_fd_sc_hd__or2_2 _29155_ (.A(_06778_),
    .B(_06645_),
    .X(_06822_));
 sky130_fd_sc_hd__a21oi_4 _29156_ (.A1(_06820_),
    .A2(_06817_),
    .B1(_06822_),
    .Y(_06823_));
 sky130_vsdinv _29157_ (.A(_06701_),
    .Y(_06824_));
 sky130_fd_sc_hd__nor2_4 _29158_ (.A(_06704_),
    .B(_06709_),
    .Y(_06825_));
 sky130_fd_sc_hd__clkbuf_4 _29159_ (.A(_19903_),
    .X(_06826_));
 sky130_fd_sc_hd__buf_6 _29160_ (.A(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__a22oi_4 _29161_ (.A1(_06502_),
    .A2(_06827_),
    .B1(_06504_),
    .B2(_06260_),
    .Y(_06828_));
 sky130_fd_sc_hd__clkbuf_2 _29162_ (.A(_06262_),
    .X(_06829_));
 sky130_fd_sc_hd__nand3_4 _29163_ (.A(_06492_),
    .B(_05404_),
    .C(_06494_),
    .Y(_06830_));
 sky130_fd_sc_hd__nor2_8 _29164_ (.A(net442),
    .B(_06830_),
    .Y(_06831_));
 sky130_fd_sc_hd__o22ai_4 _29165_ (.A1(_05261_),
    .A2(_05788_),
    .B1(_06828_),
    .B2(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2_2 _29166_ (.A(_05835_),
    .B(_19898_),
    .Y(_06833_));
 sky130_vsdinv _29167_ (.A(_06833_),
    .Y(_06834_));
 sky130_fd_sc_hd__buf_6 _29168_ (.A(_05842_),
    .X(_06835_));
 sky130_fd_sc_hd__a22o_2 _29169_ (.A1(_06502_),
    .A2(_06827_),
    .B1(_06835_),
    .B2(_05811_),
    .X(_06836_));
 sky130_fd_sc_hd__o211ai_4 _29170_ (.A1(_06272_),
    .A2(_06830_),
    .B1(_06834_),
    .C1(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__buf_6 _29171_ (.A(_06024_),
    .X(_06838_));
 sky130_fd_sc_hd__nand3_2 _29172_ (.A(_06327_),
    .B(_06838_),
    .C(_06073_),
    .Y(_06839_));
 sky130_fd_sc_hd__o22ai_4 _29173_ (.A1(net452),
    .A2(_06839_),
    .B1(_06597_),
    .B2(_06600_),
    .Y(_06840_));
 sky130_fd_sc_hd__nand3_4 _29174_ (.A(_06832_),
    .B(_06837_),
    .C(_06840_),
    .Y(_06841_));
 sky130_fd_sc_hd__o21ai_2 _29175_ (.A1(_06828_),
    .A2(_06831_),
    .B1(_06834_),
    .Y(_06842_));
 sky130_fd_sc_hd__a21oi_2 _29176_ (.A1(_06601_),
    .A2(_06598_),
    .B1(_06596_),
    .Y(_06843_));
 sky130_fd_sc_hd__o211ai_4 _29177_ (.A1(_06272_),
    .A2(_06830_),
    .B1(_06833_),
    .C1(_06836_),
    .Y(_06844_));
 sky130_fd_sc_hd__nand3_4 _29178_ (.A(_06842_),
    .B(_06843_),
    .C(_06844_),
    .Y(_06845_));
 sky130_fd_sc_hd__nor2_8 _29179_ (.A(_06691_),
    .B(_06689_),
    .Y(_06846_));
 sky130_fd_sc_hd__o2bb2ai_4 _29180_ (.A1_N(_06841_),
    .A2_N(_06845_),
    .B1(_06687_),
    .B2(_06846_),
    .Y(_06847_));
 sky130_fd_sc_hd__nor2_4 _29181_ (.A(_06687_),
    .B(_06846_),
    .Y(_06848_));
 sky130_fd_sc_hd__nand3_4 _29182_ (.A(_06845_),
    .B(_06841_),
    .C(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__o2bb2ai_4 _29183_ (.A1_N(_06623_),
    .A2_N(_06603_),
    .B1(_06614_),
    .B2(_06616_),
    .Y(_06850_));
 sky130_fd_sc_hd__a21oi_4 _29184_ (.A1(_06847_),
    .A2(_06849_),
    .B1(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__nand2_1 _29185_ (.A(_06845_),
    .B(_06848_),
    .Y(_06852_));
 sky130_vsdinv _29186_ (.A(_06841_),
    .Y(_06853_));
 sky130_fd_sc_hd__o211a_1 _29187_ (.A1(_06852_),
    .A2(_06853_),
    .B1(_06847_),
    .C1(_06850_),
    .X(_06854_));
 sky130_fd_sc_hd__o22ai_4 _29188_ (.A1(_06824_),
    .A2(_06825_),
    .B1(_06851_),
    .B2(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__and2_2 _29189_ (.A(_06710_),
    .B(_06696_),
    .X(_06856_));
 sky130_fd_sc_hd__a21o_1 _29190_ (.A1(_06847_),
    .A2(_06849_),
    .B1(_06850_),
    .X(_06857_));
 sky130_fd_sc_hd__nand3_4 _29191_ (.A(_06850_),
    .B(_06847_),
    .C(_06849_),
    .Y(_06858_));
 sky130_fd_sc_hd__nand3b_4 _29192_ (.A_N(_06856_),
    .B(_06857_),
    .C(_06858_),
    .Y(_06859_));
 sky130_vsdinv _29193_ (.A(_06717_),
    .Y(_06860_));
 sky130_fd_sc_hd__o21ai_4 _29194_ (.A1(_06860_),
    .A2(_06708_),
    .B1(_06716_),
    .Y(_06861_));
 sky130_fd_sc_hd__a21oi_4 _29195_ (.A1(_06855_),
    .A2(_06859_),
    .B1(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__a21oi_2 _29196_ (.A1(_06713_),
    .A2(_06714_),
    .B1(_06860_),
    .Y(_06863_));
 sky130_fd_sc_hd__o211a_4 _29197_ (.A1(_06711_),
    .A2(_06863_),
    .B1(_06859_),
    .C1(_06855_),
    .X(_06864_));
 sky130_fd_sc_hd__o22ai_4 _29198_ (.A1(_06821_),
    .A2(_06823_),
    .B1(_06862_),
    .B2(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__a21o_1 _29199_ (.A1(_06855_),
    .A2(_06859_),
    .B1(_06861_),
    .X(_06866_));
 sky130_fd_sc_hd__nor2_8 _29200_ (.A(_06823_),
    .B(_06821_),
    .Y(_06867_));
 sky130_fd_sc_hd__nand3_4 _29201_ (.A(_06855_),
    .B(_06861_),
    .C(_06859_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand3_4 _29202_ (.A(_06866_),
    .B(_06867_),
    .C(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand3_4 _29203_ (.A(_06865_),
    .B(_06631_),
    .C(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__o21ai_2 _29204_ (.A1(_06862_),
    .A2(_06864_),
    .B1(_06867_),
    .Y(_06871_));
 sky130_fd_sc_hd__nand3_2 _29205_ (.A(_06437_),
    .B(_06627_),
    .C(_06629_),
    .Y(_06872_));
 sky130_fd_sc_hd__a21o_1 _29206_ (.A1(_06820_),
    .A2(_06817_),
    .B1(_06822_),
    .X(_06873_));
 sky130_fd_sc_hd__nand3_1 _29207_ (.A(_06820_),
    .B(_06817_),
    .C(_06822_),
    .Y(_06874_));
 sky130_fd_sc_hd__nand2_2 _29208_ (.A(_06873_),
    .B(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__nand3_2 _29209_ (.A(_06866_),
    .B(_06868_),
    .C(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__nand3_4 _29210_ (.A(_06871_),
    .B(_06872_),
    .C(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__nor2_8 _29211_ (.A(_06729_),
    .B(_06722_),
    .Y(_06878_));
 sky130_fd_sc_hd__o2bb2ai_4 _29212_ (.A1_N(_06870_),
    .A2_N(_06877_),
    .B1(_06719_),
    .B2(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2_4 _29213_ (.A(_06730_),
    .B(_06728_),
    .Y(_06880_));
 sky130_fd_sc_hd__nand3_4 _29214_ (.A(_06877_),
    .B(_06870_),
    .C(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__clkbuf_4 _29215_ (.A(\pcpi_mul.rs2[11] ),
    .X(_06882_));
 sky130_fd_sc_hd__buf_6 _29216_ (.A(_06882_),
    .X(_06883_));
 sky130_fd_sc_hd__buf_6 _29217_ (.A(_05735_),
    .X(_06884_));
 sky130_fd_sc_hd__a22oi_4 _29218_ (.A1(_06883_),
    .A2(_05484_),
    .B1(_06884_),
    .B2(_05770_),
    .Y(_06885_));
 sky130_fd_sc_hd__nand2_1 _29219_ (.A(_06882_),
    .B(_05483_),
    .Y(_06886_));
 sky130_fd_sc_hd__nand2_1 _29220_ (.A(_06019_),
    .B(_19910_),
    .Y(_06887_));
 sky130_fd_sc_hd__nor2_1 _29221_ (.A(_06886_),
    .B(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__nand2_2 _29222_ (.A(_19659_),
    .B(_06686_),
    .Y(_06889_));
 sky130_fd_sc_hd__o21bai_1 _29223_ (.A1(_06885_),
    .A2(_06888_),
    .B1_N(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__nand3b_2 _29224_ (.A_N(_06886_),
    .B(_19655_),
    .C(_05671_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand2_1 _29225_ (.A(_06886_),
    .B(_06887_),
    .Y(_06892_));
 sky130_fd_sc_hd__nand3_1 _29226_ (.A(_06891_),
    .B(_06889_),
    .C(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__nand2_2 _29227_ (.A(_06890_),
    .B(_06893_),
    .Y(_06894_));
 sky130_vsdinv _29228_ (.A(_06894_),
    .Y(_06895_));
 sky130_fd_sc_hd__clkbuf_8 _29229_ (.A(_06605_),
    .X(_06896_));
 sky130_fd_sc_hd__buf_6 _29230_ (.A(_06167_),
    .X(_06897_));
 sky130_fd_sc_hd__buf_8 _29231_ (.A(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__a22oi_4 _29232_ (.A1(_06896_),
    .A2(_05838_),
    .B1(_06898_),
    .B2(_06330_),
    .Y(_06899_));
 sky130_fd_sc_hd__nand2_2 _29233_ (.A(_06605_),
    .B(_05695_),
    .Y(_06900_));
 sky130_fd_sc_hd__nand2_1 _29234_ (.A(_06345_),
    .B(_05236_),
    .Y(_06901_));
 sky130_fd_sc_hd__nor2_1 _29235_ (.A(_06900_),
    .B(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__nand2_2 _29236_ (.A(_06419_),
    .B(_05378_),
    .Y(_06903_));
 sky130_vsdinv _29237_ (.A(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__o21ai_1 _29238_ (.A1(_06899_),
    .A2(_06902_),
    .B1(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__buf_4 _29239_ (.A(\pcpi_mul.rs2[13] ),
    .X(_06906_));
 sky130_fd_sc_hd__buf_8 _29240_ (.A(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__nand3b_4 _29241_ (.A_N(_06900_),
    .B(_06907_),
    .C(_05225_),
    .Y(_06908_));
 sky130_fd_sc_hd__nand2_1 _29242_ (.A(_06900_),
    .B(_06901_),
    .Y(_06909_));
 sky130_fd_sc_hd__nand3_2 _29243_ (.A(_06908_),
    .B(_06903_),
    .C(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__nand2_1 _29244_ (.A(_06905_),
    .B(_06910_),
    .Y(_06911_));
 sky130_fd_sc_hd__o21ai_1 _29245_ (.A1(_06609_),
    .A2(_06611_),
    .B1(_06613_),
    .Y(_06912_));
 sky130_fd_sc_hd__and2_1 _29246_ (.A(_06912_),
    .B(_06620_),
    .X(_06913_));
 sky130_fd_sc_hd__nand2_2 _29247_ (.A(_06911_),
    .B(_06913_),
    .Y(_06914_));
 sky130_fd_sc_hd__nand2_1 _29248_ (.A(_06912_),
    .B(_06620_),
    .Y(_06915_));
 sky130_fd_sc_hd__nand3_2 _29249_ (.A(_06905_),
    .B(_06910_),
    .C(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__nand2_1 _29250_ (.A(_06914_),
    .B(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__or2_2 _29251_ (.A(_06895_),
    .B(_06917_),
    .X(_06918_));
 sky130_fd_sc_hd__nand2_2 _29252_ (.A(_06917_),
    .B(_06895_),
    .Y(_06919_));
 sky130_fd_sc_hd__buf_4 _29253_ (.A(\pcpi_mul.rs2[16] ),
    .X(_06920_));
 sky130_fd_sc_hd__clkbuf_8 _29254_ (.A(_06920_),
    .X(_06921_));
 sky130_fd_sc_hd__nand2_2 _29255_ (.A(_06921_),
    .B(_05199_),
    .Y(_06922_));
 sky130_fd_sc_hd__buf_6 _29256_ (.A(\pcpi_mul.rs2[17] ),
    .X(_06923_));
 sky130_fd_sc_hd__buf_6 _29257_ (.A(_06923_),
    .X(_06924_));
 sky130_fd_sc_hd__nand2_2 _29258_ (.A(_06924_),
    .B(_19933_),
    .Y(_06925_));
 sky130_fd_sc_hd__nor2_4 _29259_ (.A(_06922_),
    .B(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__nand2_2 _29260_ (.A(_06922_),
    .B(_06925_),
    .Y(_06927_));
 sky130_vsdinv _29261_ (.A(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__clkbuf_2 _29262_ (.A(_06433_),
    .X(_06929_));
 sky130_fd_sc_hd__nor2_4 _29263_ (.A(_06929_),
    .B(_05151_),
    .Y(_06930_));
 sky130_fd_sc_hd__o21bai_1 _29264_ (.A1(_06926_),
    .A2(_06928_),
    .B1_N(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__nand3b_1 _29265_ (.A_N(_06926_),
    .B(_06927_),
    .C(_06930_),
    .Y(_06932_));
 sky130_fd_sc_hd__nand2_2 _29266_ (.A(_06931_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__nor2_4 _29267_ (.A(_06593_),
    .B(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__and2_1 _29268_ (.A(_06933_),
    .B(_06593_),
    .X(_06935_));
 sky130_fd_sc_hd__nor2_2 _29269_ (.A(_06934_),
    .B(_06935_),
    .Y(_06936_));
 sky130_fd_sc_hd__a21o_1 _29270_ (.A1(_06918_),
    .A2(_06919_),
    .B1(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__nand3_4 _29271_ (.A(_06918_),
    .B(_06936_),
    .C(_06919_),
    .Y(_06938_));
 sky130_fd_sc_hd__nand2_1 _29272_ (.A(_06937_),
    .B(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__nand2_2 _29273_ (.A(_06939_),
    .B(_06629_),
    .Y(_06940_));
 sky130_fd_sc_hd__nand3b_4 _29274_ (.A_N(_06629_),
    .B(_06937_),
    .C(_06938_),
    .Y(_06941_));
 sky130_fd_sc_hd__nand2_4 _29275_ (.A(_06940_),
    .B(_06941_),
    .Y(_06942_));
 sky130_vsdinv _29276_ (.A(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__nand3_4 _29277_ (.A(_06879_),
    .B(_06881_),
    .C(_06943_),
    .Y(_06944_));
 sky130_vsdinv _29278_ (.A(_06941_),
    .Y(_06945_));
 sky130_vsdinv _29279_ (.A(_06940_),
    .Y(_06946_));
 sky130_fd_sc_hd__a2bb2oi_4 _29280_ (.A1_N(_06719_),
    .A2_N(_06878_),
    .B1(_06870_),
    .B2(_06877_),
    .Y(_06947_));
 sky130_fd_sc_hd__and3_1 _29281_ (.A(_06877_),
    .B(_06870_),
    .C(_06880_),
    .X(_06948_));
 sky130_fd_sc_hd__o22ai_4 _29282_ (.A1(_06945_),
    .A2(_06946_),
    .B1(_06947_),
    .B2(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__a2bb2oi_4 _29283_ (.A1_N(_06776_),
    .A2_N(_06777_),
    .B1(_06944_),
    .B2(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__a22oi_4 _29284_ (.A1(_06941_),
    .A2(_06940_),
    .B1(_06879_),
    .B2(_06881_),
    .Y(_06951_));
 sky130_fd_sc_hd__and3_1 _29285_ (.A(_06865_),
    .B(_06869_),
    .C(_06631_),
    .X(_06952_));
 sky130_fd_sc_hd__nand2_2 _29286_ (.A(_06877_),
    .B(_06880_),
    .Y(_06953_));
 sky130_fd_sc_hd__o211a_2 _29287_ (.A1(_06952_),
    .A2(_06953_),
    .B1(_06943_),
    .C1(_06879_),
    .X(_06954_));
 sky130_fd_sc_hd__nor3_4 _29288_ (.A(_06747_),
    .B(_06951_),
    .C(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__o22ai_4 _29289_ (.A1(_06774_),
    .A2(_06775_),
    .B1(_06950_),
    .B2(_06955_),
    .Y(_06956_));
 sky130_fd_sc_hd__a21boi_4 _29290_ (.A1(_06744_),
    .A2(_06589_),
    .B1_N(_06750_),
    .Y(_06957_));
 sky130_fd_sc_hd__nand2_2 _29291_ (.A(_06879_),
    .B(_06881_),
    .Y(_06958_));
 sky130_fd_sc_hd__a21oi_4 _29292_ (.A1(_06958_),
    .A2(_06942_),
    .B1(_06747_),
    .Y(_06959_));
 sky130_fd_sc_hd__nand2_2 _29293_ (.A(_06959_),
    .B(_06944_),
    .Y(_06960_));
 sky130_fd_sc_hd__o22ai_4 _29294_ (.A1(_06776_),
    .A2(_06777_),
    .B1(_06951_),
    .B2(_06954_),
    .Y(_06961_));
 sky130_fd_sc_hd__nor2_4 _29295_ (.A(_06775_),
    .B(_06774_),
    .Y(_06962_));
 sky130_fd_sc_hd__nand3_2 _29296_ (.A(_06960_),
    .B(_06961_),
    .C(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__nand3_4 _29297_ (.A(_06956_),
    .B(_06957_),
    .C(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__o21ai_2 _29298_ (.A1(_06950_),
    .A2(_06955_),
    .B1(_06962_),
    .Y(_06965_));
 sky130_vsdinv _29299_ (.A(_06957_),
    .Y(_06966_));
 sky130_vsdinv _29300_ (.A(_06962_),
    .Y(_06967_));
 sky130_fd_sc_hd__nand3_2 _29301_ (.A(_06960_),
    .B(_06961_),
    .C(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__nand3_4 _29302_ (.A(_06965_),
    .B(_06966_),
    .C(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__o2bb2ai_4 _29303_ (.A1_N(_06964_),
    .A2_N(_06969_),
    .B1(_06558_),
    .B2(_06586_),
    .Y(_06970_));
 sky130_fd_sc_hd__nand2_4 _29304_ (.A(_06964_),
    .B(_06587_),
    .Y(_06971_));
 sky130_fd_sc_hd__nand2_4 _29305_ (.A(_06768_),
    .B(_06761_),
    .Y(_06972_));
 sky130_fd_sc_hd__a21oi_4 _29306_ (.A1(_06970_),
    .A2(_06971_),
    .B1(_06972_),
    .Y(_06973_));
 sky130_fd_sc_hd__nand3_4 _29307_ (.A(_06970_),
    .B(_06972_),
    .C(_06971_),
    .Y(_06974_));
 sky130_fd_sc_hd__or2b_2 _29308_ (.A(_06973_),
    .B_N(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__o21a_1 _29309_ (.A1(_06770_),
    .A2(_06585_),
    .B1(_06769_),
    .X(_06976_));
 sky130_fd_sc_hd__xor2_4 _29310_ (.A(_06975_),
    .B(_06976_),
    .X(_02636_));
 sky130_vsdinv _29311_ (.A(_06822_),
    .Y(_06977_));
 sky130_vsdinv _29312_ (.A(_06820_),
    .Y(_06978_));
 sky130_fd_sc_hd__o21a_2 _29313_ (.A1(_06977_),
    .A2(_06978_),
    .B1(_06817_),
    .X(_06979_));
 sky130_vsdinv _29314_ (.A(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__and2_1 _29315_ (.A(_06953_),
    .B(_06870_),
    .X(_06981_));
 sky130_fd_sc_hd__nor2_2 _29316_ (.A(_06980_),
    .B(_06981_),
    .Y(_06982_));
 sky130_fd_sc_hd__nand2_4 _29317_ (.A(_06953_),
    .B(_06870_),
    .Y(_06983_));
 sky130_fd_sc_hd__nor2_2 _29318_ (.A(_06979_),
    .B(_06983_),
    .Y(_06984_));
 sky130_fd_sc_hd__nor2_2 _29319_ (.A(_06942_),
    .B(_06947_),
    .Y(_06985_));
 sky130_fd_sc_hd__buf_4 _29320_ (.A(\pcpi_mul.rs2[17] ),
    .X(_06986_));
 sky130_fd_sc_hd__nand2_2 _29321_ (.A(_06986_),
    .B(_05441_),
    .Y(_06987_));
 sky130_fd_sc_hd__buf_4 _29322_ (.A(\pcpi_mul.rs2[16] ),
    .X(_06988_));
 sky130_fd_sc_hd__nand2_2 _29323_ (.A(_06988_),
    .B(_05120_),
    .Y(_06989_));
 sky130_fd_sc_hd__nor2_4 _29324_ (.A(_06987_),
    .B(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__and2_1 _29325_ (.A(_06987_),
    .B(_06989_),
    .X(_06991_));
 sky130_fd_sc_hd__buf_4 _29326_ (.A(\pcpi_mul.rs2[15] ),
    .X(_06992_));
 sky130_fd_sc_hd__nand2_2 _29327_ (.A(_06992_),
    .B(_05467_),
    .Y(_06993_));
 sky130_vsdinv _29328_ (.A(_06993_),
    .Y(_06994_));
 sky130_fd_sc_hd__o21ai_4 _29329_ (.A1(_06990_),
    .A2(_06991_),
    .B1(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__or2_2 _29330_ (.A(_06987_),
    .B(_06989_),
    .X(_06996_));
 sky130_fd_sc_hd__nand2_2 _29331_ (.A(_06987_),
    .B(_06989_),
    .Y(_06997_));
 sky130_fd_sc_hd__nand3_4 _29332_ (.A(_06996_),
    .B(_06997_),
    .C(_06993_),
    .Y(_06998_));
 sky130_fd_sc_hd__a21oi_4 _29333_ (.A1(_06930_),
    .A2(_06927_),
    .B1(_06926_),
    .Y(_06999_));
 sky130_fd_sc_hd__nand3_4 _29334_ (.A(_06995_),
    .B(_06998_),
    .C(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__nand3_2 _29335_ (.A(_06996_),
    .B(_06997_),
    .C(_06994_),
    .Y(_07001_));
 sky130_fd_sc_hd__o21ai_2 _29336_ (.A1(_06990_),
    .A2(_06991_),
    .B1(_06993_),
    .Y(_07002_));
 sky130_fd_sc_hd__nand3b_4 _29337_ (.A_N(_06999_),
    .B(_07001_),
    .C(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__nand3_4 _29338_ (.A(_06934_),
    .B(_07000_),
    .C(_07003_),
    .Y(_07004_));
 sky130_fd_sc_hd__o2bb2ai_2 _29339_ (.A1_N(_07000_),
    .A2_N(_07003_),
    .B1(_06593_),
    .B2(_06933_),
    .Y(_07005_));
 sky130_fd_sc_hd__a22oi_4 _29340_ (.A1(_06411_),
    .A2(_05237_),
    .B1(_06343_),
    .B2(_06073_),
    .Y(_07006_));
 sky130_fd_sc_hd__buf_4 _29341_ (.A(_06413_),
    .X(_07007_));
 sky130_fd_sc_hd__buf_6 _29342_ (.A(_05172_),
    .X(_07008_));
 sky130_fd_sc_hd__nand2_2 _29343_ (.A(_07007_),
    .B(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__nand2_2 _29344_ (.A(_06897_),
    .B(_05271_),
    .Y(_07010_));
 sky130_fd_sc_hd__nor2_2 _29345_ (.A(_07009_),
    .B(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__nand2_2 _29346_ (.A(_19649_),
    .B(_05486_),
    .Y(_07012_));
 sky130_fd_sc_hd__o21ai_2 _29347_ (.A1(_07006_),
    .A2(_07011_),
    .B1(_07012_),
    .Y(_07013_));
 sky130_fd_sc_hd__nand3b_2 _29348_ (.A_N(_07009_),
    .B(_06618_),
    .C(_19918_),
    .Y(_07014_));
 sky130_vsdinv _29349_ (.A(_07012_),
    .Y(_07015_));
 sky130_fd_sc_hd__nand2_2 _29350_ (.A(_07009_),
    .B(_07010_),
    .Y(_07016_));
 sky130_fd_sc_hd__nand3_2 _29351_ (.A(_07014_),
    .B(_07015_),
    .C(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__o21ai_2 _29352_ (.A1(_06903_),
    .A2(_06899_),
    .B1(_06908_),
    .Y(_07018_));
 sky130_fd_sc_hd__nand3_4 _29353_ (.A(_07013_),
    .B(_07017_),
    .C(_07018_),
    .Y(_07019_));
 sky130_fd_sc_hd__o21ai_2 _29354_ (.A1(_07006_),
    .A2(_07011_),
    .B1(_07015_),
    .Y(_07020_));
 sky130_fd_sc_hd__nand3_2 _29355_ (.A(_07014_),
    .B(_07012_),
    .C(_07016_),
    .Y(_07021_));
 sky130_fd_sc_hd__o21ai_1 _29356_ (.A1(_06900_),
    .A2(_06901_),
    .B1(_06903_),
    .Y(_07022_));
 sky130_fd_sc_hd__nand2_1 _29357_ (.A(_07022_),
    .B(_06909_),
    .Y(_07023_));
 sky130_fd_sc_hd__nand3_4 _29358_ (.A(_07020_),
    .B(_07021_),
    .C(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__a22oi_4 _29359_ (.A1(net477),
    .A2(_05666_),
    .B1(_19655_),
    .B2(_06106_),
    .Y(_07025_));
 sky130_fd_sc_hd__nand2_1 _29360_ (.A(_06401_),
    .B(_05481_),
    .Y(_07026_));
 sky130_fd_sc_hd__nand2_1 _29361_ (.A(_19654_),
    .B(_05672_),
    .Y(_07027_));
 sky130_fd_sc_hd__nor2_2 _29362_ (.A(_07026_),
    .B(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__nand2_2 _29363_ (.A(_06013_),
    .B(_05673_),
    .Y(_07029_));
 sky130_fd_sc_hd__o21bai_2 _29364_ (.A1(_07025_),
    .A2(_07028_),
    .B1_N(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__nand3b_2 _29365_ (.A_N(_07026_),
    .B(_06838_),
    .C(_05808_),
    .Y(_07031_));
 sky130_fd_sc_hd__nand2_1 _29366_ (.A(_07026_),
    .B(_07027_),
    .Y(_07032_));
 sky130_fd_sc_hd__nand3_2 _29367_ (.A(_07031_),
    .B(_07032_),
    .C(_07029_),
    .Y(_07033_));
 sky130_fd_sc_hd__nand2_4 _29368_ (.A(_07030_),
    .B(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__a21o_1 _29369_ (.A1(_07019_),
    .A2(_07024_),
    .B1(_07034_),
    .X(_07035_));
 sky130_fd_sc_hd__nand3_2 _29370_ (.A(_07019_),
    .B(_07024_),
    .C(_07034_),
    .Y(_07036_));
 sky130_fd_sc_hd__nand2_2 _29371_ (.A(_07035_),
    .B(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__a21o_1 _29372_ (.A1(_07004_),
    .A2(_07005_),
    .B1(_07037_),
    .X(_07038_));
 sky130_fd_sc_hd__nand3_4 _29373_ (.A(_07037_),
    .B(_07004_),
    .C(_07005_),
    .Y(_07039_));
 sky130_fd_sc_hd__a21o_2 _29374_ (.A1(_07038_),
    .A2(_07039_),
    .B1(_06938_),
    .X(_07040_));
 sky130_fd_sc_hd__clkinv_8 _29375_ (.A(\pcpi_mul.rs2[18] ),
    .Y(_07041_));
 sky130_fd_sc_hd__buf_4 _29376_ (.A(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__nor2_4 _29377_ (.A(_07042_),
    .B(_04842_),
    .Y(_07043_));
 sky130_fd_sc_hd__nand3_4 _29378_ (.A(_06938_),
    .B(_07038_),
    .C(_07039_),
    .Y(_07044_));
 sky130_fd_sc_hd__and3_4 _29379_ (.A(_07040_),
    .B(_07043_),
    .C(_07044_),
    .X(_07045_));
 sky130_fd_sc_hd__a21oi_4 _29380_ (.A1(_07040_),
    .A2(_07044_),
    .B1(_07043_),
    .Y(_07046_));
 sky130_fd_sc_hd__nor2_8 _29381_ (.A(_06867_),
    .B(_06864_),
    .Y(_07047_));
 sky130_fd_sc_hd__nor2_4 _29382_ (.A(_06802_),
    .B(_06800_),
    .Y(_07048_));
 sky130_fd_sc_hd__a21bo_1 _29383_ (.A1(_06793_),
    .A2(_06812_),
    .B1_N(_06797_),
    .X(_07049_));
 sky130_fd_sc_hd__buf_4 _29384_ (.A(\pcpi_mul.rs1[17] ),
    .X(_07050_));
 sky130_fd_sc_hd__buf_6 _29385_ (.A(_07050_),
    .X(_07051_));
 sky130_fd_sc_hd__buf_6 _29386_ (.A(_06798_),
    .X(_07052_));
 sky130_fd_sc_hd__nand2_1 _29387_ (.A(_06636_),
    .B(_07052_),
    .Y(_07053_));
 sky130_fd_sc_hd__a21o_1 _29388_ (.A1(_05223_),
    .A2(_07051_),
    .B1(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__buf_6 _29389_ (.A(_19880_),
    .X(_07055_));
 sky130_fd_sc_hd__buf_6 _29390_ (.A(_07050_),
    .X(_07056_));
 sky130_fd_sc_hd__nand2_1 _29391_ (.A(_05163_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__a21o_1 _29392_ (.A1(_06639_),
    .A2(_07055_),
    .B1(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__buf_6 _29393_ (.A(_19883_),
    .X(_07059_));
 sky130_fd_sc_hd__buf_6 _29394_ (.A(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__nand2_2 _29395_ (.A(_05157_),
    .B(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__nand3_2 _29396_ (.A(_07054_),
    .B(_07058_),
    .C(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__a21o_1 _29397_ (.A1(_07054_),
    .A2(_07058_),
    .B1(_07061_),
    .X(_07063_));
 sky130_fd_sc_hd__buf_4 _29398_ (.A(_06808_),
    .X(_07064_));
 sky130_fd_sc_hd__a22oi_4 _29399_ (.A1(_05768_),
    .A2(_19891_),
    .B1(_05647_),
    .B2(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__and4_1 _29400_ (.A(_05778_),
    .B(_05169_),
    .C(_19888_),
    .D(_06462_),
    .X(_07066_));
 sky130_fd_sc_hd__clkbuf_8 _29401_ (.A(\pcpi_mul.rs1[18] ),
    .X(_07067_));
 sky130_fd_sc_hd__nand2_4 _29402_ (.A(_05290_),
    .B(_07067_),
    .Y(_07068_));
 sky130_vsdinv _29403_ (.A(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__o21ai_2 _29404_ (.A1(_07065_),
    .A2(_07066_),
    .B1(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__a21oi_2 _29405_ (.A1(_06791_),
    .A2(_06785_),
    .B1(_06782_),
    .Y(_07071_));
 sky130_fd_sc_hd__buf_6 _29406_ (.A(_06282_),
    .X(_07072_));
 sky130_fd_sc_hd__nand2_1 _29407_ (.A(_05772_),
    .B(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__nand3b_4 _29408_ (.A_N(_07073_),
    .B(_06659_),
    .C(_06640_),
    .Y(_07074_));
 sky130_fd_sc_hd__a22o_1 _29409_ (.A1(_05212_),
    .A2(_19891_),
    .B1(_05647_),
    .B2(_07064_),
    .X(_07075_));
 sky130_fd_sc_hd__nand3_2 _29410_ (.A(_07074_),
    .B(_07075_),
    .C(_07068_),
    .Y(_07076_));
 sky130_fd_sc_hd__nand3_4 _29411_ (.A(_07070_),
    .B(_07071_),
    .C(_07076_),
    .Y(_07077_));
 sky130_fd_sc_hd__o21ai_2 _29412_ (.A1(_07065_),
    .A2(_07066_),
    .B1(_07068_),
    .Y(_07078_));
 sky130_fd_sc_hd__nand3_4 _29413_ (.A(_07074_),
    .B(_07075_),
    .C(_07069_),
    .Y(_07079_));
 sky130_fd_sc_hd__o21ai_4 _29414_ (.A1(_06784_),
    .A2(_06781_),
    .B1(_06790_),
    .Y(_07080_));
 sky130_fd_sc_hd__nand3_4 _29415_ (.A(_07078_),
    .B(_07079_),
    .C(_07080_),
    .Y(_07081_));
 sky130_fd_sc_hd__a22o_2 _29416_ (.A1(_07062_),
    .A2(_07063_),
    .B1(_07077_),
    .B2(_07081_),
    .X(_07082_));
 sky130_fd_sc_hd__a21oi_2 _29417_ (.A1(_07054_),
    .A2(_07058_),
    .B1(_07061_),
    .Y(_07083_));
 sky130_fd_sc_hd__and3_1 _29418_ (.A(_07054_),
    .B(_07058_),
    .C(_07061_),
    .X(_07084_));
 sky130_fd_sc_hd__nor2_4 _29419_ (.A(_07083_),
    .B(_07084_),
    .Y(_07085_));
 sky130_fd_sc_hd__nand3_4 _29420_ (.A(_07085_),
    .B(_07077_),
    .C(_07081_),
    .Y(_07086_));
 sky130_fd_sc_hd__nand3_4 _29421_ (.A(_07049_),
    .B(_07082_),
    .C(_07086_),
    .Y(_07087_));
 sky130_vsdinv _29422_ (.A(_06793_),
    .Y(_07088_));
 sky130_fd_sc_hd__o21a_1 _29423_ (.A1(_06811_),
    .A2(_06807_),
    .B1(_06797_),
    .X(_07089_));
 sky130_fd_sc_hd__o2bb2ai_4 _29424_ (.A1_N(_07086_),
    .A2_N(_07082_),
    .B1(_07088_),
    .B2(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__o211a_1 _29425_ (.A1(_07048_),
    .A2(_06807_),
    .B1(_07087_),
    .C1(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__or2_2 _29426_ (.A(_07048_),
    .B(_06807_),
    .X(_07092_));
 sky130_fd_sc_hd__a21oi_4 _29427_ (.A1(_07090_),
    .A2(_07087_),
    .B1(_07092_),
    .Y(_07093_));
 sky130_fd_sc_hd__nand2_1 _29428_ (.A(_06858_),
    .B(_06856_),
    .Y(_07094_));
 sky130_vsdinv _29429_ (.A(_06845_),
    .Y(_07095_));
 sky130_fd_sc_hd__nor2_2 _29430_ (.A(_06848_),
    .B(_06853_),
    .Y(_07096_));
 sky130_fd_sc_hd__a22oi_4 _29431_ (.A1(_05451_),
    .A2(_19901_),
    .B1(_05833_),
    .B2(_05774_),
    .Y(_07097_));
 sky130_fd_sc_hd__nand3_4 _29432_ (.A(_05586_),
    .B(_05842_),
    .C(_05798_),
    .Y(_07098_));
 sky130_fd_sc_hd__nor2_8 _29433_ (.A(_05787_),
    .B(_07098_),
    .Y(_07099_));
 sky130_fd_sc_hd__o22ai_4 _29434_ (.A1(_05261_),
    .A2(_06471_),
    .B1(_07097_),
    .B2(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__o21ai_2 _29435_ (.A1(_06889_),
    .A2(_06885_),
    .B1(_06891_),
    .Y(_07101_));
 sky130_fd_sc_hd__buf_6 _29436_ (.A(_05787_),
    .X(_07102_));
 sky130_fd_sc_hd__nand2_2 _29437_ (.A(_19667_),
    .B(_06288_),
    .Y(_07103_));
 sky130_vsdinv _29438_ (.A(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__a22o_2 _29439_ (.A1(_05832_),
    .A2(_05804_),
    .B1(_06488_),
    .B2(_06649_),
    .X(_07105_));
 sky130_fd_sc_hd__o211ai_4 _29440_ (.A1(_07102_),
    .A2(_07098_),
    .B1(_07104_),
    .C1(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__nand3_4 _29441_ (.A(_07100_),
    .B(_07101_),
    .C(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__o21ai_2 _29442_ (.A1(_07097_),
    .A2(_07099_),
    .B1(_07104_),
    .Y(_07108_));
 sky130_fd_sc_hd__o21ai_1 _29443_ (.A1(_06886_),
    .A2(_06887_),
    .B1(_06889_),
    .Y(_07109_));
 sky130_fd_sc_hd__nand2_1 _29444_ (.A(_07109_),
    .B(_06892_),
    .Y(_07110_));
 sky130_fd_sc_hd__o211ai_4 _29445_ (.A1(_05788_),
    .A2(_07098_),
    .B1(_07103_),
    .C1(_07105_),
    .Y(_07111_));
 sky130_fd_sc_hd__nand3_4 _29446_ (.A(_07108_),
    .B(_07110_),
    .C(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__nor2_8 _29447_ (.A(_06834_),
    .B(_06831_),
    .Y(_07113_));
 sky130_fd_sc_hd__o2bb2ai_4 _29448_ (.A1_N(_07107_),
    .A2_N(_07112_),
    .B1(_06828_),
    .B2(_07113_),
    .Y(_07114_));
 sky130_fd_sc_hd__nor2_4 _29449_ (.A(_06828_),
    .B(_07113_),
    .Y(_07115_));
 sky130_fd_sc_hd__nand3_4 _29450_ (.A(_07112_),
    .B(_07107_),
    .C(_07115_),
    .Y(_07116_));
 sky130_fd_sc_hd__nand2_2 _29451_ (.A(_06916_),
    .B(_06894_),
    .Y(_07117_));
 sky130_fd_sc_hd__nand2_4 _29452_ (.A(_07117_),
    .B(_06914_),
    .Y(_07118_));
 sky130_fd_sc_hd__a21oi_4 _29453_ (.A1(_07114_),
    .A2(_07116_),
    .B1(_07118_),
    .Y(_07119_));
 sky130_vsdinv _29454_ (.A(_07107_),
    .Y(_07120_));
 sky130_fd_sc_hd__nand2_1 _29455_ (.A(_07112_),
    .B(_07115_),
    .Y(_07121_));
 sky130_fd_sc_hd__o211a_1 _29456_ (.A1(_07120_),
    .A2(_07121_),
    .B1(_07114_),
    .C1(_07118_),
    .X(_07122_));
 sky130_fd_sc_hd__o22ai_4 _29457_ (.A1(_07095_),
    .A2(_07096_),
    .B1(_07119_),
    .B2(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__nand2_1 _29458_ (.A(_07114_),
    .B(_07116_),
    .Y(_07124_));
 sky130_fd_sc_hd__and2_1 _29459_ (.A(_07117_),
    .B(_06914_),
    .X(_07125_));
 sky130_fd_sc_hd__nand2_2 _29460_ (.A(_07124_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__nand3_4 _29461_ (.A(_07118_),
    .B(_07114_),
    .C(_07116_),
    .Y(_07127_));
 sky130_fd_sc_hd__nand2_2 _29462_ (.A(_06852_),
    .B(_06841_),
    .Y(_07128_));
 sky130_fd_sc_hd__nand3_4 _29463_ (.A(_07126_),
    .B(_07127_),
    .C(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__a22oi_4 _29464_ (.A1(_06857_),
    .A2(_07094_),
    .B1(_07123_),
    .B2(_07129_),
    .Y(_07130_));
 sky130_vsdinv _29465_ (.A(_06849_),
    .Y(_07131_));
 sky130_fd_sc_hd__o2bb2ai_1 _29466_ (.A1_N(_07125_),
    .A2_N(_07124_),
    .B1(_06853_),
    .B2(_07131_),
    .Y(_07132_));
 sky130_fd_sc_hd__o21ai_4 _29467_ (.A1(_06856_),
    .A2(_06851_),
    .B1(_06858_),
    .Y(_07133_));
 sky130_fd_sc_hd__o211a_2 _29468_ (.A1(_07122_),
    .A2(_07132_),
    .B1(_07133_),
    .C1(_07123_),
    .X(_07134_));
 sky130_fd_sc_hd__o22ai_4 _29469_ (.A1(_07091_),
    .A2(_07093_),
    .B1(_07130_),
    .B2(_07134_),
    .Y(_07135_));
 sky130_fd_sc_hd__a21o_1 _29470_ (.A1(_07123_),
    .A2(_07129_),
    .B1(_07133_),
    .X(_07136_));
 sky130_fd_sc_hd__nor2_2 _29471_ (.A(_07093_),
    .B(_07091_),
    .Y(_07137_));
 sky130_fd_sc_hd__nand3_4 _29472_ (.A(_07123_),
    .B(_07133_),
    .C(_07129_),
    .Y(_07138_));
 sky130_fd_sc_hd__nand3_2 _29473_ (.A(_07136_),
    .B(_07137_),
    .C(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__nand3_1 _29474_ (.A(_07135_),
    .B(_06945_),
    .C(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__clkbuf_4 _29475_ (.A(_07140_),
    .X(_07141_));
 sky130_fd_sc_hd__o21ai_2 _29476_ (.A1(_07130_),
    .A2(_07134_),
    .B1(_07137_),
    .Y(_07142_));
 sky130_fd_sc_hd__a21o_1 _29477_ (.A1(_07090_),
    .A2(_07087_),
    .B1(_07092_),
    .X(_07143_));
 sky130_fd_sc_hd__nand3_1 _29478_ (.A(_07090_),
    .B(_07092_),
    .C(_07087_),
    .Y(_07144_));
 sky130_fd_sc_hd__nand2_2 _29479_ (.A(_07143_),
    .B(_07144_),
    .Y(_07145_));
 sky130_fd_sc_hd__nand3_2 _29480_ (.A(_07136_),
    .B(_07138_),
    .C(_07145_),
    .Y(_07146_));
 sky130_fd_sc_hd__nand3_4 _29481_ (.A(_07142_),
    .B(_06941_),
    .C(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__a2bb2oi_2 _29482_ (.A1_N(_06862_),
    .A2_N(_07047_),
    .B1(_07141_),
    .B2(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__nor2_2 _29483_ (.A(_06862_),
    .B(_06875_),
    .Y(_07149_));
 sky130_fd_sc_hd__o211a_1 _29484_ (.A1(_06864_),
    .A2(_07149_),
    .B1(_07140_),
    .C1(_07147_),
    .X(_07150_));
 sky130_fd_sc_hd__o22ai_4 _29485_ (.A1(_07045_),
    .A2(_07046_),
    .B1(_07148_),
    .B2(_07150_),
    .Y(_07151_));
 sky130_fd_sc_hd__o2bb2ai_4 _29486_ (.A1_N(_07141_),
    .A2_N(_07147_),
    .B1(_06862_),
    .B2(_07047_),
    .Y(_07152_));
 sky130_fd_sc_hd__nor2_8 _29487_ (.A(_07046_),
    .B(_07045_),
    .Y(_07153_));
 sky130_fd_sc_hd__nor2_4 _29488_ (.A(_06862_),
    .B(_07047_),
    .Y(_07154_));
 sky130_fd_sc_hd__nand3_4 _29489_ (.A(_07147_),
    .B(_07154_),
    .C(_07141_),
    .Y(_07155_));
 sky130_fd_sc_hd__nand3_4 _29490_ (.A(_07152_),
    .B(_07153_),
    .C(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__a22oi_4 _29491_ (.A1(_06985_),
    .A2(_06881_),
    .B1(_07151_),
    .B2(_07156_),
    .Y(_07157_));
 sky130_fd_sc_hd__nand2_1 _29492_ (.A(_07147_),
    .B(_07141_),
    .Y(_07158_));
 sky130_fd_sc_hd__nor2_2 _29493_ (.A(_06864_),
    .B(_07149_),
    .Y(_07159_));
 sky130_fd_sc_hd__a21boi_4 _29494_ (.A1(_07158_),
    .A2(_07159_),
    .B1_N(_07153_),
    .Y(_07160_));
 sky130_fd_sc_hd__a21oi_4 _29495_ (.A1(_07152_),
    .A2(_07155_),
    .B1(_07153_),
    .Y(_07161_));
 sky130_fd_sc_hd__a211oi_4 _29496_ (.A1(_07155_),
    .A2(_07160_),
    .B1(_06944_),
    .C1(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__o22ai_4 _29497_ (.A1(_06982_),
    .A2(_06984_),
    .B1(_07157_),
    .B2(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__a22oi_4 _29498_ (.A1(_06944_),
    .A2(_06959_),
    .B1(_06961_),
    .B2(_06967_),
    .Y(_07164_));
 sky130_fd_sc_hd__and3_1 _29499_ (.A(_07135_),
    .B(_07139_),
    .C(_06945_),
    .X(_07165_));
 sky130_fd_sc_hd__nand2_2 _29500_ (.A(_07147_),
    .B(_07154_),
    .Y(_07166_));
 sky130_fd_sc_hd__o211a_4 _29501_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07153_),
    .C1(_07152_),
    .X(_07167_));
 sky130_fd_sc_hd__nand2_2 _29502_ (.A(_06954_),
    .B(_07151_),
    .Y(_07168_));
 sky130_fd_sc_hd__nand2_1 _29503_ (.A(_06981_),
    .B(_06979_),
    .Y(_07169_));
 sky130_fd_sc_hd__nand2_4 _29504_ (.A(_06983_),
    .B(_06980_),
    .Y(_07170_));
 sky130_fd_sc_hd__nand2_4 _29505_ (.A(_07169_),
    .B(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__o22ai_4 _29506_ (.A1(_06942_),
    .A2(_06958_),
    .B1(_07161_),
    .B2(_07167_),
    .Y(_07172_));
 sky130_fd_sc_hd__o211ai_4 _29507_ (.A1(_07167_),
    .A2(_07168_),
    .B1(_07171_),
    .C1(_07172_),
    .Y(_07173_));
 sky130_fd_sc_hd__nand3_4 _29508_ (.A(_07163_),
    .B(_07164_),
    .C(_07173_),
    .Y(_07174_));
 sky130_fd_sc_hd__xor2_2 _29509_ (.A(_06980_),
    .B(_06983_),
    .X(_07175_));
 sky130_fd_sc_hd__nand2_1 _29510_ (.A(_07172_),
    .B(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__o21ai_2 _29511_ (.A1(_06962_),
    .A2(_06950_),
    .B1(_06960_),
    .Y(_07177_));
 sky130_fd_sc_hd__o21ai_2 _29512_ (.A1(_07157_),
    .A2(_07162_),
    .B1(_07171_),
    .Y(_07178_));
 sky130_fd_sc_hd__o211ai_4 _29513_ (.A1(_07162_),
    .A2(_07176_),
    .B1(_07177_),
    .C1(_07178_),
    .Y(_07179_));
 sky130_vsdinv _29514_ (.A(_06773_),
    .Y(_07180_));
 sky130_fd_sc_hd__o2bb2ai_2 _29515_ (.A1_N(_07174_),
    .A2_N(_07179_),
    .B1(_06732_),
    .B2(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__nor2_4 _29516_ (.A(_07180_),
    .B(_06732_),
    .Y(_07182_));
 sky130_fd_sc_hd__nand2_8 _29517_ (.A(_07174_),
    .B(_07182_),
    .Y(_07183_));
 sky130_fd_sc_hd__nand2_2 _29518_ (.A(_06971_),
    .B(_06969_),
    .Y(_07184_));
 sky130_fd_sc_hd__a21oi_4 _29519_ (.A1(_07181_),
    .A2(_07183_),
    .B1(_07184_),
    .Y(_07185_));
 sky130_vsdinv _29520_ (.A(_07185_),
    .Y(_07186_));
 sky130_fd_sc_hd__nand2_2 _29521_ (.A(_06970_),
    .B(_06971_),
    .Y(_07187_));
 sky130_vsdinv _29522_ (.A(_06972_),
    .Y(_07188_));
 sky130_fd_sc_hd__a21oi_4 _29523_ (.A1(_07187_),
    .A2(_07188_),
    .B1(_06770_),
    .Y(_07189_));
 sky130_fd_sc_hd__a21oi_4 _29524_ (.A1(_06769_),
    .A2(_06974_),
    .B1(_06973_),
    .Y(_07190_));
 sky130_fd_sc_hd__a31o_2 _29525_ (.A1(_06584_),
    .A2(_06974_),
    .A3(_07189_),
    .B1(_07190_),
    .X(_07191_));
 sky130_fd_sc_hd__nand2_1 _29526_ (.A(_07179_),
    .B(_07174_),
    .Y(_07192_));
 sky130_vsdinv _29527_ (.A(_07182_),
    .Y(_07193_));
 sky130_fd_sc_hd__a22oi_4 _29528_ (.A1(_06971_),
    .A2(_06969_),
    .B1(_07192_),
    .B2(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__a21oi_4 _29529_ (.A1(_07183_),
    .A2(_07194_),
    .B1(_07185_),
    .Y(_07195_));
 sky130_fd_sc_hd__nor2_2 _29530_ (.A(_07195_),
    .B(_07191_),
    .Y(_07196_));
 sky130_fd_sc_hd__a21oi_4 _29531_ (.A1(_07186_),
    .A2(_07191_),
    .B1(_07196_),
    .Y(_02637_));
 sky130_fd_sc_hd__a21oi_2 _29532_ (.A1(_07172_),
    .A2(_07175_),
    .B1(_07162_),
    .Y(_07197_));
 sky130_fd_sc_hd__a21oi_4 _29533_ (.A1(_06995_),
    .A2(_06998_),
    .B1(_06999_),
    .Y(_07198_));
 sky130_fd_sc_hd__a21o_1 _29534_ (.A1(_06994_),
    .A2(_06997_),
    .B1(_06990_),
    .X(_07199_));
 sky130_fd_sc_hd__inv_4 _29535_ (.A(_19919_),
    .Y(_07200_));
 sky130_fd_sc_hd__nor2_4 _29536_ (.A(_06433_),
    .B(_07200_),
    .Y(_07201_));
 sky130_vsdinv _29537_ (.A(_07201_),
    .Y(_07202_));
 sky130_fd_sc_hd__nand2_2 _29538_ (.A(_06923_),
    .B(_05229_),
    .Y(_07203_));
 sky130_fd_sc_hd__nand2_2 _29539_ (.A(_06920_),
    .B(_19923_),
    .Y(_07204_));
 sky130_fd_sc_hd__nor2_4 _29540_ (.A(_07203_),
    .B(_07204_),
    .Y(_07205_));
 sky130_vsdinv _29541_ (.A(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__nand2_2 _29542_ (.A(_07203_),
    .B(_07204_),
    .Y(_07207_));
 sky130_fd_sc_hd__nand3_2 _29543_ (.A(_07202_),
    .B(_07206_),
    .C(_07207_),
    .Y(_07208_));
 sky130_vsdinv _29544_ (.A(_07207_),
    .Y(_07209_));
 sky130_fd_sc_hd__o21ai_2 _29545_ (.A1(_07205_),
    .A2(_07209_),
    .B1(_07201_),
    .Y(_07210_));
 sky130_fd_sc_hd__nand3b_4 _29546_ (.A_N(_07199_),
    .B(_07208_),
    .C(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__o21ai_2 _29547_ (.A1(_07205_),
    .A2(_07209_),
    .B1(_07202_),
    .Y(_07212_));
 sky130_fd_sc_hd__nand3_2 _29548_ (.A(_07206_),
    .B(_07207_),
    .C(_07201_),
    .Y(_07213_));
 sky130_fd_sc_hd__nand3_4 _29549_ (.A(_07212_),
    .B(_07213_),
    .C(_07199_),
    .Y(_07214_));
 sky130_fd_sc_hd__nand3_4 _29550_ (.A(_07198_),
    .B(_07211_),
    .C(_07214_),
    .Y(_07215_));
 sky130_fd_sc_hd__a21o_1 _29551_ (.A1(_07211_),
    .A2(_07214_),
    .B1(_07198_),
    .X(_07216_));
 sky130_fd_sc_hd__o21ai_1 _29552_ (.A1(_07009_),
    .A2(_07010_),
    .B1(_07012_),
    .Y(_07217_));
 sky130_fd_sc_hd__and2_1 _29553_ (.A(_07217_),
    .B(_07016_),
    .X(_07218_));
 sky130_fd_sc_hd__a22oi_4 _29554_ (.A1(_06414_),
    .A2(_05268_),
    .B1(_06345_),
    .B2(_05637_),
    .Y(_07219_));
 sky130_fd_sc_hd__nand2_2 _29555_ (.A(_06413_),
    .B(_05267_),
    .Y(_07220_));
 sky130_fd_sc_hd__nand2_2 _29556_ (.A(_06897_),
    .B(_05379_),
    .Y(_07221_));
 sky130_fd_sc_hd__nor2_2 _29557_ (.A(_07220_),
    .B(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__buf_4 _29558_ (.A(\pcpi_mul.rs2[12] ),
    .X(_07223_));
 sky130_fd_sc_hd__nand2_2 _29559_ (.A(_07223_),
    .B(_05769_),
    .Y(_07224_));
 sky130_fd_sc_hd__o21ai_2 _29560_ (.A1(_07219_),
    .A2(_07222_),
    .B1(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__nand3b_4 _29561_ (.A_N(_07220_),
    .B(_06416_),
    .C(_05380_),
    .Y(_07226_));
 sky130_vsdinv _29562_ (.A(_07224_),
    .Y(_07227_));
 sky130_fd_sc_hd__nand2_2 _29563_ (.A(_07220_),
    .B(_07221_),
    .Y(_07228_));
 sky130_fd_sc_hd__nand3_2 _29564_ (.A(_07226_),
    .B(_07227_),
    .C(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__nand3_4 _29565_ (.A(_07218_),
    .B(_07225_),
    .C(_07229_),
    .Y(_07230_));
 sky130_fd_sc_hd__o21ai_2 _29566_ (.A1(_07219_),
    .A2(_07222_),
    .B1(_07227_),
    .Y(_07231_));
 sky130_fd_sc_hd__nand3_2 _29567_ (.A(_07226_),
    .B(_07224_),
    .C(_07228_),
    .Y(_07232_));
 sky130_fd_sc_hd__nand2_1 _29568_ (.A(_07217_),
    .B(_07016_),
    .Y(_07233_));
 sky130_fd_sc_hd__nand3_4 _29569_ (.A(_07231_),
    .B(_07232_),
    .C(_07233_),
    .Y(_07234_));
 sky130_fd_sc_hd__a22oi_4 _29570_ (.A1(_06022_),
    .A2(_05661_),
    .B1(_05736_),
    .B2(_06494_),
    .Y(_07235_));
 sky130_fd_sc_hd__nand2_1 _29571_ (.A(_06017_),
    .B(_05463_),
    .Y(_07236_));
 sky130_fd_sc_hd__nand2_1 _29572_ (.A(_06158_),
    .B(_06826_),
    .Y(_07237_));
 sky130_fd_sc_hd__nor2_1 _29573_ (.A(_07236_),
    .B(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__nand2_2 _29574_ (.A(_06013_),
    .B(_05798_),
    .Y(_07239_));
 sky130_fd_sc_hd__o21bai_2 _29575_ (.A1(_07235_),
    .A2(_07238_),
    .B1_N(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__nand3b_2 _29576_ (.A_N(_07236_),
    .B(_06884_),
    .C(_06257_),
    .Y(_07241_));
 sky130_fd_sc_hd__nand2_1 _29577_ (.A(_07236_),
    .B(_07237_),
    .Y(_07242_));
 sky130_fd_sc_hd__nand3_2 _29578_ (.A(_07241_),
    .B(_07239_),
    .C(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__nand2_4 _29579_ (.A(_07240_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__a21oi_1 _29580_ (.A1(_07230_),
    .A2(_07234_),
    .B1(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__nand2_2 _29581_ (.A(_07234_),
    .B(_07244_),
    .Y(_07246_));
 sky130_vsdinv _29582_ (.A(_07230_),
    .Y(_07247_));
 sky130_fd_sc_hd__nor2_1 _29583_ (.A(_07246_),
    .B(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__o2bb2ai_2 _29584_ (.A1_N(_07215_),
    .A2_N(_07216_),
    .B1(_07245_),
    .B2(_07248_),
    .Y(_07249_));
 sky130_fd_sc_hd__nand3_1 _29585_ (.A(_07005_),
    .B(_07036_),
    .C(_07035_),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_1 _29586_ (.A(_07250_),
    .B(_07004_),
    .Y(_07251_));
 sky130_fd_sc_hd__a21o_1 _29587_ (.A1(_07230_),
    .A2(_07234_),
    .B1(_07244_),
    .X(_07252_));
 sky130_fd_sc_hd__o2111ai_4 _29588_ (.A1(_07246_),
    .A2(_07247_),
    .B1(_07215_),
    .C1(_07252_),
    .D1(_07216_),
    .Y(_07253_));
 sky130_fd_sc_hd__nand3_4 _29589_ (.A(_07249_),
    .B(_07251_),
    .C(_07253_),
    .Y(_07254_));
 sky130_fd_sc_hd__nand2_1 _29590_ (.A(_07249_),
    .B(_07253_),
    .Y(_07255_));
 sky130_fd_sc_hd__and2_1 _29591_ (.A(_07250_),
    .B(_07004_),
    .X(_07256_));
 sky130_fd_sc_hd__nand2_2 _29592_ (.A(_07255_),
    .B(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__buf_4 _29593_ (.A(\pcpi_mul.rs2[19] ),
    .X(_07258_));
 sky130_fd_sc_hd__nand2_2 _29594_ (.A(_07258_),
    .B(\pcpi_mul.rs1[0] ),
    .Y(_07259_));
 sky130_fd_sc_hd__nand2_4 _29595_ (.A(\pcpi_mul.rs2[18] ),
    .B(_19929_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_1 _29596_ (.A(_07259_),
    .B(_07260_),
    .Y(_07261_));
 sky130_vsdinv _29597_ (.A(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__nor2_4 _29598_ (.A(_07259_),
    .B(_07260_),
    .Y(_07263_));
 sky130_fd_sc_hd__o2bb2ai_2 _29599_ (.A1_N(_07254_),
    .A2_N(_07257_),
    .B1(_07262_),
    .B2(_07263_),
    .Y(_07264_));
 sky130_vsdinv _29600_ (.A(_07263_),
    .Y(_07265_));
 sky130_fd_sc_hd__nand2_1 _29601_ (.A(_07265_),
    .B(_07261_),
    .Y(_07266_));
 sky130_vsdinv _29602_ (.A(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__nand3_4 _29603_ (.A(_07257_),
    .B(_07254_),
    .C(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__nand3_2 _29604_ (.A(_07040_),
    .B(_07043_),
    .C(_07044_),
    .Y(_07269_));
 sky130_fd_sc_hd__a21boi_4 _29605_ (.A1(_07264_),
    .A2(_07268_),
    .B1_N(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__clkbuf_4 _29606_ (.A(_07268_),
    .X(_07271_));
 sky130_fd_sc_hd__and3_1 _29607_ (.A(_07045_),
    .B(_07264_),
    .C(_07271_),
    .X(_07272_));
 sky130_vsdinv _29608_ (.A(_07121_),
    .Y(_07273_));
 sky130_vsdinv _29609_ (.A(_06282_),
    .Y(_07274_));
 sky130_fd_sc_hd__buf_6 _29610_ (.A(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__a22oi_4 _29611_ (.A1(_05446_),
    .A2(_06440_),
    .B1(_05447_),
    .B2(_06652_),
    .Y(_07276_));
 sky130_fd_sc_hd__nand3_4 _29612_ (.A(_05586_),
    .B(_05588_),
    .C(_06118_),
    .Y(_07277_));
 sky130_fd_sc_hd__nor2_8 _29613_ (.A(_06460_),
    .B(_07277_),
    .Y(_07278_));
 sky130_fd_sc_hd__o22ai_4 _29614_ (.A1(_05261_),
    .A2(_07275_),
    .B1(_07276_),
    .B2(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__o21ai_2 _29615_ (.A1(_07029_),
    .A2(_07025_),
    .B1(_07031_),
    .Y(_07280_));
 sky130_fd_sc_hd__buf_6 _29616_ (.A(_06282_),
    .X(_07281_));
 sky130_fd_sc_hd__and2_4 _29617_ (.A(_05699_),
    .B(_07281_),
    .X(_07282_));
 sky130_fd_sc_hd__a22o_2 _29618_ (.A1(_05446_),
    .A2(_06440_),
    .B1(_06217_),
    .B2(_19894_),
    .X(_07283_));
 sky130_fd_sc_hd__o211ai_4 _29619_ (.A1(_06471_),
    .A2(_07277_),
    .B1(_07282_),
    .C1(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__nand3_4 _29620_ (.A(_07279_),
    .B(_07280_),
    .C(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__o21ai_2 _29621_ (.A1(_07276_),
    .A2(_07278_),
    .B1(_07282_),
    .Y(_07286_));
 sky130_vsdinv _29622_ (.A(_07029_),
    .Y(_07287_));
 sky130_fd_sc_hd__a21oi_2 _29623_ (.A1(_07287_),
    .A2(_07032_),
    .B1(_07028_),
    .Y(_07288_));
 sky130_fd_sc_hd__clkbuf_2 _29624_ (.A(_07274_),
    .X(_07289_));
 sky130_fd_sc_hd__o221ai_4 _29625_ (.A1(_05260_),
    .A2(_07289_),
    .B1(_06460_),
    .B2(_07277_),
    .C1(_07283_),
    .Y(_07290_));
 sky130_fd_sc_hd__nand3_4 _29626_ (.A(_07286_),
    .B(_07288_),
    .C(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__nor2_8 _29627_ (.A(_07104_),
    .B(_07099_),
    .Y(_07292_));
 sky130_fd_sc_hd__o2bb2ai_4 _29628_ (.A1_N(_07285_),
    .A2_N(_07291_),
    .B1(_07097_),
    .B2(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__nor2_2 _29629_ (.A(_07097_),
    .B(_07292_),
    .Y(_07294_));
 sky130_fd_sc_hd__nand3_4 _29630_ (.A(_07291_),
    .B(_07285_),
    .C(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__nand2_1 _29631_ (.A(_07024_),
    .B(_07034_),
    .Y(_07296_));
 sky130_fd_sc_hd__nand2_4 _29632_ (.A(_07296_),
    .B(_07019_),
    .Y(_07297_));
 sky130_fd_sc_hd__a21oi_4 _29633_ (.A1(_07293_),
    .A2(_07295_),
    .B1(_07297_),
    .Y(_07298_));
 sky130_vsdinv _29634_ (.A(_07285_),
    .Y(_07299_));
 sky130_fd_sc_hd__nand2_1 _29635_ (.A(_07291_),
    .B(_07294_),
    .Y(_07300_));
 sky130_fd_sc_hd__o211a_2 _29636_ (.A1(_07299_),
    .A2(_07300_),
    .B1(_07293_),
    .C1(_07297_),
    .X(_07301_));
 sky130_fd_sc_hd__o22ai_4 _29637_ (.A1(_07120_),
    .A2(_07273_),
    .B1(_07298_),
    .B2(_07301_),
    .Y(_07302_));
 sky130_vsdinv _29638_ (.A(_07128_),
    .Y(_07303_));
 sky130_fd_sc_hd__nand2_1 _29639_ (.A(_07127_),
    .B(_07303_),
    .Y(_07304_));
 sky130_fd_sc_hd__nand2_1 _29640_ (.A(_07304_),
    .B(_07126_),
    .Y(_07305_));
 sky130_fd_sc_hd__a21o_1 _29641_ (.A1(_07293_),
    .A2(_07295_),
    .B1(_07297_),
    .X(_07306_));
 sky130_fd_sc_hd__nand3_4 _29642_ (.A(_07297_),
    .B(_07293_),
    .C(_07295_),
    .Y(_07307_));
 sky130_fd_sc_hd__nor2_4 _29643_ (.A(_07120_),
    .B(_07273_),
    .Y(_07308_));
 sky130_fd_sc_hd__nand3_2 _29644_ (.A(_07306_),
    .B(_07307_),
    .C(_07308_),
    .Y(_07309_));
 sky130_fd_sc_hd__nand3_4 _29645_ (.A(_07302_),
    .B(_07305_),
    .C(_07309_),
    .Y(_07310_));
 sky130_vsdinv _29646_ (.A(_07112_),
    .Y(_07311_));
 sky130_fd_sc_hd__nor2_2 _29647_ (.A(_07115_),
    .B(_07120_),
    .Y(_07312_));
 sky130_fd_sc_hd__o22ai_4 _29648_ (.A1(_07311_),
    .A2(_07312_),
    .B1(_07298_),
    .B2(_07301_),
    .Y(_07313_));
 sky130_fd_sc_hd__o21ai_2 _29649_ (.A1(_07303_),
    .A2(_07119_),
    .B1(_07127_),
    .Y(_07314_));
 sky130_fd_sc_hd__o211ai_2 _29650_ (.A1(_07120_),
    .A2(_07273_),
    .B1(_07307_),
    .C1(_07306_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand3_4 _29651_ (.A(_07313_),
    .B(_07314_),
    .C(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__nand2_1 _29652_ (.A(_07310_),
    .B(_07316_),
    .Y(_07317_));
 sky130_fd_sc_hd__a21oi_2 _29653_ (.A1(_07078_),
    .A2(_07079_),
    .B1(_07080_),
    .Y(_07318_));
 sky130_fd_sc_hd__nand2_1 _29654_ (.A(_07063_),
    .B(_07062_),
    .Y(_07319_));
 sky130_fd_sc_hd__o21ai_4 _29655_ (.A1(_07318_),
    .A2(_07319_),
    .B1(_07081_),
    .Y(_07320_));
 sky130_fd_sc_hd__nand2_1 _29656_ (.A(_05280_),
    .B(_06464_),
    .Y(_07321_));
 sky130_fd_sc_hd__buf_6 _29657_ (.A(\pcpi_mul.rs1[15] ),
    .X(_07322_));
 sky130_fd_sc_hd__buf_6 _29658_ (.A(_07322_),
    .X(_07323_));
 sky130_fd_sc_hd__nand3b_4 _29659_ (.A_N(_07321_),
    .B(_06659_),
    .C(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__buf_6 _29660_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07325_));
 sky130_fd_sc_hd__nand2_4 _29661_ (.A(_05171_),
    .B(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__buf_6 _29662_ (.A(_19887_),
    .X(_07327_));
 sky130_fd_sc_hd__a22o_1 _29663_ (.A1(_05212_),
    .A2(_07327_),
    .B1(_05792_),
    .B2(_06635_),
    .X(_07328_));
 sky130_fd_sc_hd__nand3_2 _29664_ (.A(_07324_),
    .B(_07326_),
    .C(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__buf_6 _29665_ (.A(_19886_),
    .X(_07330_));
 sky130_fd_sc_hd__a22oi_4 _29666_ (.A1(_05295_),
    .A2(_07330_),
    .B1(_19673_),
    .B2(_19884_),
    .Y(_07331_));
 sky130_fd_sc_hd__and4_2 _29667_ (.A(_05768_),
    .B(_06258_),
    .C(_06641_),
    .D(_19888_),
    .X(_07332_));
 sky130_vsdinv _29668_ (.A(_07326_),
    .Y(_07333_));
 sky130_fd_sc_hd__o21ai_2 _29669_ (.A1(_07331_),
    .A2(_07332_),
    .B1(_07333_),
    .Y(_07334_));
 sky130_fd_sc_hd__o2111ai_4 _29670_ (.A1(_07065_),
    .A2(_07068_),
    .B1(_07074_),
    .C1(_07329_),
    .D1(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__o21ai_4 _29671_ (.A1(_07331_),
    .A2(_07332_),
    .B1(_07326_),
    .Y(_07336_));
 sky130_fd_sc_hd__nand3_4 _29672_ (.A(_07324_),
    .B(_07333_),
    .C(_07328_),
    .Y(_07337_));
 sky130_fd_sc_hd__o21ai_4 _29673_ (.A1(_07068_),
    .A2(_07065_),
    .B1(_07074_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand3_4 _29674_ (.A(_07336_),
    .B(_07337_),
    .C(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__nand2_1 _29675_ (.A(_07335_),
    .B(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand2_2 _29676_ (.A(_06639_),
    .B(_19878_),
    .Y(_07341_));
 sky130_fd_sc_hd__a21o_2 _29677_ (.A1(_05164_),
    .A2(_19874_),
    .B1(_07341_),
    .X(_07342_));
 sky130_fd_sc_hd__clkbuf_8 _29678_ (.A(\pcpi_mul.rs1[17] ),
    .X(_07343_));
 sky130_fd_sc_hd__buf_6 _29679_ (.A(_07343_),
    .X(_07344_));
 sky130_fd_sc_hd__buf_4 _29680_ (.A(\pcpi_mul.rs1[18] ),
    .X(_07345_));
 sky130_fd_sc_hd__buf_6 _29681_ (.A(_07345_),
    .X(_07346_));
 sky130_fd_sc_hd__nand2_2 _29682_ (.A(_19683_),
    .B(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__a21o_2 _29683_ (.A1(_05162_),
    .A2(_07344_),
    .B1(_07347_),
    .X(_07348_));
 sky130_fd_sc_hd__nand2_4 _29684_ (.A(_19677_),
    .B(net454),
    .Y(_07349_));
 sky130_fd_sc_hd__a21o_1 _29685_ (.A1(_07342_),
    .A2(_07348_),
    .B1(_07349_),
    .X(_07350_));
 sky130_fd_sc_hd__nand3_4 _29686_ (.A(_07342_),
    .B(_07348_),
    .C(_07349_),
    .Y(_07351_));
 sky130_fd_sc_hd__nand2_4 _29687_ (.A(_07350_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__nand2_1 _29688_ (.A(_07340_),
    .B(_07352_),
    .Y(_07353_));
 sky130_fd_sc_hd__a21oi_4 _29689_ (.A1(_07342_),
    .A2(_07348_),
    .B1(_07349_),
    .Y(_07354_));
 sky130_vsdinv _29690_ (.A(_07351_),
    .Y(_07355_));
 sky130_fd_sc_hd__nor2_2 _29691_ (.A(_07354_),
    .B(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__nand3_2 _29692_ (.A(_07356_),
    .B(_07335_),
    .C(_07339_),
    .Y(_07357_));
 sky130_fd_sc_hd__nand3_4 _29693_ (.A(_07320_),
    .B(_07353_),
    .C(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__a21boi_4 _29694_ (.A1(_07085_),
    .A2(_07077_),
    .B1_N(_07081_),
    .Y(_07359_));
 sky130_fd_sc_hd__nand2_2 _29695_ (.A(_07340_),
    .B(_07356_),
    .Y(_07360_));
 sky130_fd_sc_hd__nand3_4 _29696_ (.A(_07352_),
    .B(_07335_),
    .C(_07339_),
    .Y(_07361_));
 sky130_fd_sc_hd__o21a_4 _29697_ (.A1(_07053_),
    .A2(_07057_),
    .B1(_07063_),
    .X(_07362_));
 sky130_fd_sc_hd__a31oi_4 _29698_ (.A1(_07359_),
    .A2(_07360_),
    .A3(_07361_),
    .B1(_07362_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand3_4 _29699_ (.A(_07359_),
    .B(_07360_),
    .C(_07361_),
    .Y(_07364_));
 sky130_fd_sc_hd__a21boi_4 _29700_ (.A1(_07364_),
    .A2(_07358_),
    .B1_N(_07362_),
    .Y(_07365_));
 sky130_fd_sc_hd__a21oi_2 _29701_ (.A1(_07358_),
    .A2(_07363_),
    .B1(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__nand2_1 _29702_ (.A(_07317_),
    .B(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__nand2_1 _29703_ (.A(_07364_),
    .B(_07358_),
    .Y(_07368_));
 sky130_fd_sc_hd__nor2_4 _29704_ (.A(_07362_),
    .B(_07368_),
    .Y(_07369_));
 sky130_fd_sc_hd__o211ai_4 _29705_ (.A1(_07365_),
    .A2(_07369_),
    .B1(_07310_),
    .C1(_07316_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand3_4 _29706_ (.A(_07367_),
    .B(_07040_),
    .C(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__o2bb2ai_2 _29707_ (.A1_N(_07316_),
    .A2_N(_07310_),
    .B1(_07369_),
    .B2(_07365_),
    .Y(_07372_));
 sky130_vsdinv _29708_ (.A(_07040_),
    .Y(_07373_));
 sky130_fd_sc_hd__nand3_2 _29709_ (.A(_07366_),
    .B(_07310_),
    .C(_07316_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand3_4 _29710_ (.A(_07372_),
    .B(_07373_),
    .C(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__o21ai_4 _29711_ (.A1(_07130_),
    .A2(_07145_),
    .B1(_07138_),
    .Y(_07376_));
 sky130_fd_sc_hd__a21oi_2 _29712_ (.A1(_07371_),
    .A2(_07375_),
    .B1(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__nor2_1 _29713_ (.A(_07130_),
    .B(_07145_),
    .Y(_07378_));
 sky130_fd_sc_hd__o211a_1 _29714_ (.A1(_07134_),
    .A2(_07378_),
    .B1(_07375_),
    .C1(_07371_),
    .X(_07379_));
 sky130_fd_sc_hd__o22ai_4 _29715_ (.A1(_07270_),
    .A2(_07272_),
    .B1(_07377_),
    .B2(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__a21o_1 _29716_ (.A1(_07371_),
    .A2(_07375_),
    .B1(_07376_),
    .X(_07381_));
 sky130_fd_sc_hd__nand2_1 _29717_ (.A(_07257_),
    .B(_07254_),
    .Y(_07382_));
 sky130_fd_sc_hd__a21oi_1 _29718_ (.A1(_07382_),
    .A2(_07266_),
    .B1(_07269_),
    .Y(_07383_));
 sky130_fd_sc_hd__a21oi_2 _29719_ (.A1(_07271_),
    .A2(_07383_),
    .B1(_07270_),
    .Y(_07384_));
 sky130_fd_sc_hd__nand3_4 _29720_ (.A(_07371_),
    .B(_07375_),
    .C(_07376_),
    .Y(_07385_));
 sky130_fd_sc_hd__nand3_4 _29721_ (.A(_07381_),
    .B(_07384_),
    .C(_07385_),
    .Y(_07386_));
 sky130_fd_sc_hd__a21boi_4 _29722_ (.A1(_07380_),
    .A2(_07386_),
    .B1_N(_07156_),
    .Y(_07387_));
 sky130_fd_sc_hd__o2111a_1 _29723_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07160_),
    .C1(_07386_),
    .D1(_07380_),
    .X(_07388_));
 sky130_fd_sc_hd__nand2_2 _29724_ (.A(_07166_),
    .B(_07141_),
    .Y(_07389_));
 sky130_vsdinv _29725_ (.A(_07092_),
    .Y(_07390_));
 sky130_vsdinv _29726_ (.A(_07090_),
    .Y(_07391_));
 sky130_fd_sc_hd__o21a_2 _29727_ (.A1(_07390_),
    .A2(_07391_),
    .B1(_07087_),
    .X(_07392_));
 sky130_vsdinv _29728_ (.A(_07392_),
    .Y(_07393_));
 sky130_fd_sc_hd__nand2_4 _29729_ (.A(_07389_),
    .B(_07393_),
    .Y(_07394_));
 sky130_fd_sc_hd__nand3_2 _29730_ (.A(_07166_),
    .B(_07141_),
    .C(_07392_),
    .Y(_07395_));
 sky130_fd_sc_hd__nand2_4 _29731_ (.A(_07394_),
    .B(_07395_),
    .Y(_07396_));
 sky130_fd_sc_hd__o21bai_2 _29732_ (.A1(_07387_),
    .A2(_07388_),
    .B1_N(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__a21o_1 _29733_ (.A1(_07386_),
    .A2(_07380_),
    .B1(_07167_),
    .X(_07398_));
 sky130_fd_sc_hd__nand3_4 _29734_ (.A(_07167_),
    .B(_07386_),
    .C(_07380_),
    .Y(_07399_));
 sky130_fd_sc_hd__nand3_2 _29735_ (.A(_07398_),
    .B(_07396_),
    .C(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__nand3_4 _29736_ (.A(_07197_),
    .B(_07397_),
    .C(_07400_),
    .Y(_07401_));
 sky130_fd_sc_hd__o21ai_2 _29737_ (.A1(_07387_),
    .A2(_07388_),
    .B1(_07396_),
    .Y(_07402_));
 sky130_fd_sc_hd__o22ai_4 _29738_ (.A1(_07167_),
    .A2(_07168_),
    .B1(_07171_),
    .B2(_07157_),
    .Y(_07403_));
 sky130_vsdinv _29739_ (.A(_07396_),
    .Y(_07404_));
 sky130_fd_sc_hd__nand3_2 _29740_ (.A(_07398_),
    .B(_07404_),
    .C(_07399_),
    .Y(_07405_));
 sky130_fd_sc_hd__nand3_4 _29741_ (.A(_07402_),
    .B(_07403_),
    .C(_07405_),
    .Y(_07406_));
 sky130_fd_sc_hd__nand2_1 _29742_ (.A(_07401_),
    .B(_07406_),
    .Y(_07407_));
 sky130_fd_sc_hd__a22oi_4 _29743_ (.A1(_07407_),
    .A2(_07170_),
    .B1(_07179_),
    .B2(_07183_),
    .Y(_07408_));
 sky130_vsdinv _29744_ (.A(_07170_),
    .Y(_07409_));
 sky130_fd_sc_hd__nand3_4 _29745_ (.A(_07401_),
    .B(_07406_),
    .C(_07409_),
    .Y(_07410_));
 sky130_fd_sc_hd__o2bb2ai_2 _29746_ (.A1_N(_07406_),
    .A2_N(_07401_),
    .B1(_06979_),
    .B2(_06981_),
    .Y(_07411_));
 sky130_fd_sc_hd__nand2_1 _29747_ (.A(_07183_),
    .B(_07179_),
    .Y(_07412_));
 sky130_fd_sc_hd__a21oi_4 _29748_ (.A1(_07411_),
    .A2(_07410_),
    .B1(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__a21oi_4 _29749_ (.A1(_07408_),
    .A2(_07410_),
    .B1(_07413_),
    .Y(_07414_));
 sky130_fd_sc_hd__a22oi_4 _29750_ (.A1(_07183_),
    .A2(_07194_),
    .B1(_07191_),
    .B2(_07195_),
    .Y(_07415_));
 sky130_fd_sc_hd__xnor2_4 _29751_ (.A(_07414_),
    .B(_07415_),
    .Y(_02638_));
 sky130_fd_sc_hd__nor2b_4 _29752_ (.A(_07363_),
    .B_N(_07358_),
    .Y(_07416_));
 sky130_fd_sc_hd__nand2_2 _29753_ (.A(_07385_),
    .B(_07375_),
    .Y(_07417_));
 sky130_vsdinv _29754_ (.A(_07417_),
    .Y(_07418_));
 sky130_fd_sc_hd__nor2_8 _29755_ (.A(_07416_),
    .B(_07418_),
    .Y(_07419_));
 sky130_fd_sc_hd__and3_1 _29756_ (.A(_07385_),
    .B(_07375_),
    .C(_07416_),
    .X(_07420_));
 sky130_fd_sc_hd__a22oi_4 _29757_ (.A1(_19631_),
    .A2(_05146_),
    .B1(_19635_),
    .B2(_05236_),
    .Y(_07421_));
 sky130_fd_sc_hd__nand3_4 _29758_ (.A(_06923_),
    .B(_06920_),
    .C(_05263_),
    .Y(_07422_));
 sky130_fd_sc_hd__nor2_4 _29759_ (.A(_07200_),
    .B(_07422_),
    .Y(_07423_));
 sky130_fd_sc_hd__nand2_2 _29760_ (.A(_06992_),
    .B(_05271_),
    .Y(_07424_));
 sky130_fd_sc_hd__o21ai_2 _29761_ (.A1(_07421_),
    .A2(_07423_),
    .B1(_07424_),
    .Y(_07425_));
 sky130_fd_sc_hd__buf_6 _29762_ (.A(_07200_),
    .X(_07426_));
 sky130_vsdinv _29763_ (.A(_07424_),
    .Y(_07427_));
 sky130_fd_sc_hd__buf_6 _29764_ (.A(\pcpi_mul.rs2[16] ),
    .X(_07428_));
 sky130_fd_sc_hd__a22o_2 _29765_ (.A1(_06986_),
    .A2(_05467_),
    .B1(_07428_),
    .B2(_07008_),
    .X(_07429_));
 sky130_fd_sc_hd__o211ai_4 _29766_ (.A1(_07426_),
    .A2(_07422_),
    .B1(_07427_),
    .C1(_07429_),
    .Y(_07430_));
 sky130_fd_sc_hd__nand3_4 _29767_ (.A(_07425_),
    .B(_07263_),
    .C(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__o21ai_2 _29768_ (.A1(_07421_),
    .A2(_07423_),
    .B1(_07427_),
    .Y(_07432_));
 sky130_fd_sc_hd__o211ai_4 _29769_ (.A1(_07200_),
    .A2(_07422_),
    .B1(_07424_),
    .C1(_07429_),
    .Y(_07433_));
 sky130_fd_sc_hd__nand3_4 _29770_ (.A(_07432_),
    .B(_07265_),
    .C(_07433_),
    .Y(_07434_));
 sky130_fd_sc_hd__buf_6 _29771_ (.A(_06992_),
    .X(_07435_));
 sky130_fd_sc_hd__a31o_2 _29772_ (.A1(_07207_),
    .A2(_07435_),
    .A3(_19921_),
    .B1(_07205_),
    .X(_07436_));
 sky130_fd_sc_hd__a21o_1 _29773_ (.A1(_07431_),
    .A2(_07434_),
    .B1(_07436_),
    .X(_07437_));
 sky130_vsdinv _29774_ (.A(_07214_),
    .Y(_07438_));
 sky130_fd_sc_hd__nand3_4 _29775_ (.A(_07431_),
    .B(_07434_),
    .C(_07436_),
    .Y(_07439_));
 sky130_fd_sc_hd__nand3_4 _29776_ (.A(_07437_),
    .B(_07438_),
    .C(_07439_),
    .Y(_07440_));
 sky130_fd_sc_hd__a21oi_2 _29777_ (.A1(_07431_),
    .A2(_07434_),
    .B1(_07436_),
    .Y(_07441_));
 sky130_fd_sc_hd__and3_1 _29778_ (.A(_07431_),
    .B(_07434_),
    .C(_07436_),
    .X(_07442_));
 sky130_fd_sc_hd__o21ai_4 _29779_ (.A1(_07441_),
    .A2(_07442_),
    .B1(_07214_),
    .Y(_07443_));
 sky130_fd_sc_hd__a22oi_4 _29780_ (.A1(_19644_),
    .A2(_05380_),
    .B1(_06422_),
    .B2(_05489_),
    .Y(_07444_));
 sky130_fd_sc_hd__nand2_2 _29781_ (.A(_19643_),
    .B(_05379_),
    .Y(_07445_));
 sky130_fd_sc_hd__nand2_2 _29782_ (.A(_19646_),
    .B(_05488_),
    .Y(_07446_));
 sky130_fd_sc_hd__nor2_4 _29783_ (.A(_07445_),
    .B(_07446_),
    .Y(_07447_));
 sky130_fd_sc_hd__nand2_2 _29784_ (.A(\pcpi_mul.rs2[12] ),
    .B(_05660_),
    .Y(_07448_));
 sky130_fd_sc_hd__o21ai_2 _29785_ (.A1(_07444_),
    .A2(_07447_),
    .B1(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__nand3b_4 _29786_ (.A_N(_07445_),
    .B(_06907_),
    .C(_05666_),
    .Y(_07450_));
 sky130_vsdinv _29787_ (.A(_07448_),
    .Y(_07451_));
 sky130_fd_sc_hd__nand2_4 _29788_ (.A(_07445_),
    .B(_07446_),
    .Y(_07452_));
 sky130_fd_sc_hd__nand3_4 _29789_ (.A(_07450_),
    .B(_07451_),
    .C(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__o21ai_2 _29790_ (.A1(_07224_),
    .A2(_07219_),
    .B1(_07226_),
    .Y(_07454_));
 sky130_fd_sc_hd__nand3_4 _29791_ (.A(_07449_),
    .B(_07453_),
    .C(_07454_),
    .Y(_07455_));
 sky130_fd_sc_hd__o21ai_2 _29792_ (.A1(_07444_),
    .A2(_07447_),
    .B1(_07451_),
    .Y(_07456_));
 sky130_fd_sc_hd__nand3_2 _29793_ (.A(_07450_),
    .B(_07448_),
    .C(_07452_),
    .Y(_07457_));
 sky130_fd_sc_hd__o21ai_1 _29794_ (.A1(_07220_),
    .A2(_07221_),
    .B1(_07224_),
    .Y(_07458_));
 sky130_fd_sc_hd__nand2_1 _29795_ (.A(_07458_),
    .B(_07228_),
    .Y(_07459_));
 sky130_fd_sc_hd__nand3_4 _29796_ (.A(_07456_),
    .B(_07457_),
    .C(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__a22oi_4 _29797_ (.A1(_06018_),
    .A2(_06494_),
    .B1(_06019_),
    .B2(_05804_),
    .Y(_07461_));
 sky130_fd_sc_hd__nand2_1 _29798_ (.A(_06882_),
    .B(_05558_),
    .Y(_07462_));
 sky130_fd_sc_hd__nand2_1 _29799_ (.A(_05882_),
    .B(_05798_),
    .Y(_07463_));
 sky130_fd_sc_hd__nor2_2 _29800_ (.A(_07462_),
    .B(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__nand2_2 _29801_ (.A(_19658_),
    .B(_06118_),
    .Y(_07465_));
 sky130_vsdinv _29802_ (.A(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__o21ai_2 _29803_ (.A1(_07461_),
    .A2(_07464_),
    .B1(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__nand3b_4 _29804_ (.A_N(_07462_),
    .B(_06884_),
    .C(_05811_),
    .Y(_07468_));
 sky130_fd_sc_hd__nand2_1 _29805_ (.A(_07462_),
    .B(_07463_),
    .Y(_07469_));
 sky130_fd_sc_hd__nand3_2 _29806_ (.A(_07468_),
    .B(_07465_),
    .C(_07469_),
    .Y(_07470_));
 sky130_fd_sc_hd__nand2_4 _29807_ (.A(_07467_),
    .B(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__nand3_1 _29808_ (.A(_07455_),
    .B(_07460_),
    .C(_07471_),
    .Y(_07472_));
 sky130_vsdinv _29809_ (.A(_07472_),
    .Y(_07473_));
 sky130_fd_sc_hd__a21oi_4 _29810_ (.A1(_07455_),
    .A2(_07460_),
    .B1(_07471_),
    .Y(_07474_));
 sky130_fd_sc_hd__o2bb2ai_4 _29811_ (.A1_N(_07440_),
    .A2_N(_07443_),
    .B1(_07473_),
    .B2(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__nor2_4 _29812_ (.A(_07474_),
    .B(_07473_),
    .Y(_07476_));
 sky130_fd_sc_hd__nand3_4 _29813_ (.A(_07443_),
    .B(_07476_),
    .C(_07440_),
    .Y(_07477_));
 sky130_fd_sc_hd__nand2_2 _29814_ (.A(_07253_),
    .B(_07215_),
    .Y(_07478_));
 sky130_fd_sc_hd__a21oi_2 _29815_ (.A1(_07475_),
    .A2(_07477_),
    .B1(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__and3_2 _29816_ (.A(_07475_),
    .B(_07478_),
    .C(_07477_),
    .X(_07480_));
 sky130_fd_sc_hd__buf_4 _29817_ (.A(\pcpi_mul.rs2[18] ),
    .X(_07481_));
 sky130_fd_sc_hd__nand2_2 _29818_ (.A(_07481_),
    .B(_19927_),
    .Y(_07482_));
 sky130_fd_sc_hd__nand2_1 _29819_ (.A(_07258_),
    .B(_05105_),
    .Y(_07483_));
 sky130_fd_sc_hd__buf_6 _29820_ (.A(_19621_),
    .X(_07484_));
 sky130_fd_sc_hd__nand3b_2 _29821_ (.A_N(_07483_),
    .B(_07484_),
    .C(_05213_),
    .Y(_07485_));
 sky130_fd_sc_hd__buf_4 _29822_ (.A(_19620_),
    .X(_07486_));
 sky130_fd_sc_hd__nand2_1 _29823_ (.A(_07486_),
    .B(_05198_),
    .Y(_07487_));
 sky130_fd_sc_hd__nand2_1 _29824_ (.A(_07483_),
    .B(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__and2_1 _29825_ (.A(_07485_),
    .B(_07488_),
    .X(_07489_));
 sky130_fd_sc_hd__or2_1 _29826_ (.A(_07482_),
    .B(_07489_),
    .X(_07490_));
 sky130_fd_sc_hd__nand2_1 _29827_ (.A(_07489_),
    .B(_07482_),
    .Y(_07491_));
 sky130_fd_sc_hd__nand2_2 _29828_ (.A(_07490_),
    .B(_07491_),
    .Y(_07492_));
 sky130_vsdinv _29829_ (.A(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__o21ai_4 _29830_ (.A1(_07479_),
    .A2(_07480_),
    .B1(_07493_),
    .Y(_07494_));
 sky130_fd_sc_hd__a21o_1 _29831_ (.A1(_07475_),
    .A2(_07477_),
    .B1(_07478_),
    .X(_07495_));
 sky130_fd_sc_hd__nand3_4 _29832_ (.A(_07475_),
    .B(_07478_),
    .C(_07477_),
    .Y(_07496_));
 sky130_fd_sc_hd__nand3_4 _29833_ (.A(_07495_),
    .B(_07496_),
    .C(_07492_),
    .Y(_07497_));
 sky130_fd_sc_hd__a21boi_4 _29834_ (.A1(_07494_),
    .A2(_07497_),
    .B1_N(_07271_),
    .Y(_07498_));
 sky130_fd_sc_hd__nand2_2 _29835_ (.A(_07494_),
    .B(_07497_),
    .Y(_07499_));
 sky130_fd_sc_hd__nor2_2 _29836_ (.A(_07271_),
    .B(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__a22oi_4 _29837_ (.A1(_05451_),
    .A2(_06788_),
    .B1(_06488_),
    .B2(_06462_),
    .Y(_07501_));
 sky130_fd_sc_hd__buf_6 _29838_ (.A(_06287_),
    .X(_07502_));
 sky130_fd_sc_hd__nand3_4 _29839_ (.A(_05586_),
    .B(_05588_),
    .C(_07502_),
    .Y(_07503_));
 sky130_fd_sc_hd__nor2_8 _29840_ (.A(_07274_),
    .B(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__nand2_2 _29841_ (.A(_05443_),
    .B(_06267_),
    .Y(_07505_));
 sky130_fd_sc_hd__o21ai_2 _29842_ (.A1(_07501_),
    .A2(_07504_),
    .B1(_07505_),
    .Y(_07506_));
 sky130_fd_sc_hd__o21ai_2 _29843_ (.A1(_07239_),
    .A2(_07235_),
    .B1(_07241_),
    .Y(_07507_));
 sky130_vsdinv _29844_ (.A(_07505_),
    .Y(_07508_));
 sky130_fd_sc_hd__a22o_1 _29845_ (.A1(_19662_),
    .A2(_05962_),
    .B1(_06488_),
    .B2(_07281_),
    .X(_07509_));
 sky130_fd_sc_hd__o211ai_2 _29846_ (.A1(_07275_),
    .A2(_07503_),
    .B1(_07508_),
    .C1(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__nand3_4 _29847_ (.A(_07506_),
    .B(_07507_),
    .C(_07510_),
    .Y(_07511_));
 sky130_fd_sc_hd__o21ai_2 _29848_ (.A1(_07501_),
    .A2(_07504_),
    .B1(_07508_),
    .Y(_07512_));
 sky130_fd_sc_hd__o21ai_1 _29849_ (.A1(_07236_),
    .A2(_07237_),
    .B1(_07239_),
    .Y(_07513_));
 sky130_fd_sc_hd__nand2_1 _29850_ (.A(_07513_),
    .B(_07242_),
    .Y(_07514_));
 sky130_fd_sc_hd__o211ai_2 _29851_ (.A1(_07275_),
    .A2(_07503_),
    .B1(_07505_),
    .C1(_07509_),
    .Y(_07515_));
 sky130_fd_sc_hd__nand3_4 _29852_ (.A(_07512_),
    .B(_07514_),
    .C(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__nor2_8 _29853_ (.A(_07282_),
    .B(_07278_),
    .Y(_07517_));
 sky130_fd_sc_hd__o2bb2ai_4 _29854_ (.A1_N(_07511_),
    .A2_N(_07516_),
    .B1(_07276_),
    .B2(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__nor2_2 _29855_ (.A(_07276_),
    .B(_07517_),
    .Y(_07519_));
 sky130_fd_sc_hd__nand3_4 _29856_ (.A(_07511_),
    .B(_07516_),
    .C(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__nand2_4 _29857_ (.A(_07246_),
    .B(_07230_),
    .Y(_07521_));
 sky130_fd_sc_hd__a21oi_4 _29858_ (.A1(_07518_),
    .A2(_07520_),
    .B1(_07521_),
    .Y(_07522_));
 sky130_fd_sc_hd__nand2_1 _29859_ (.A(_07516_),
    .B(_07519_),
    .Y(_07523_));
 sky130_vsdinv _29860_ (.A(_07511_),
    .Y(_07524_));
 sky130_fd_sc_hd__o211a_1 _29861_ (.A1(_07523_),
    .A2(_07524_),
    .B1(_07518_),
    .C1(_07521_),
    .X(_07525_));
 sky130_fd_sc_hd__nand2_2 _29862_ (.A(_07300_),
    .B(_07285_),
    .Y(_07526_));
 sky130_vsdinv _29863_ (.A(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__o21ai_4 _29864_ (.A1(_07522_),
    .A2(_07525_),
    .B1(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__a21o_1 _29865_ (.A1(_07518_),
    .A2(_07520_),
    .B1(_07521_),
    .X(_07529_));
 sky130_fd_sc_hd__nand3_4 _29866_ (.A(_07521_),
    .B(_07518_),
    .C(_07520_),
    .Y(_07530_));
 sky130_fd_sc_hd__nand3_4 _29867_ (.A(_07529_),
    .B(_07530_),
    .C(_07526_),
    .Y(_07531_));
 sky130_fd_sc_hd__o21ai_4 _29868_ (.A1(_07308_),
    .A2(_07298_),
    .B1(_07307_),
    .Y(_07532_));
 sky130_fd_sc_hd__a21oi_4 _29869_ (.A1(_07528_),
    .A2(_07531_),
    .B1(_07532_),
    .Y(_07533_));
 sky130_fd_sc_hd__nor2_1 _29870_ (.A(_07308_),
    .B(_07298_),
    .Y(_07534_));
 sky130_fd_sc_hd__o211a_2 _29871_ (.A1(_07301_),
    .A2(_07534_),
    .B1(_07531_),
    .C1(_07528_),
    .X(_07535_));
 sky130_fd_sc_hd__nor2_4 _29872_ (.A(_07341_),
    .B(_07347_),
    .Y(_07536_));
 sky130_fd_sc_hd__a21oi_4 _29873_ (.A1(_07336_),
    .A2(_07337_),
    .B1(_07338_),
    .Y(_07537_));
 sky130_fd_sc_hd__o21ai_4 _29874_ (.A1(_07326_),
    .A2(_07331_),
    .B1(_07324_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand2_4 _29875_ (.A(_05211_),
    .B(_07322_),
    .Y(_07539_));
 sky130_fd_sc_hd__nand2_4 _29876_ (.A(_05201_),
    .B(_19880_),
    .Y(_07540_));
 sky130_fd_sc_hd__or2_2 _29877_ (.A(_07539_),
    .B(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__buf_6 _29878_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07542_));
 sky130_fd_sc_hd__nand2_4 _29879_ (.A(_19685_),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__nand2_4 _29880_ (.A(_07539_),
    .B(_07540_),
    .Y(_07544_));
 sky130_fd_sc_hd__nand3_2 _29881_ (.A(_07541_),
    .B(_07543_),
    .C(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__a22oi_4 _29882_ (.A1(_05768_),
    .A2(_06641_),
    .B1(_05647_),
    .B2(_07052_),
    .Y(_07546_));
 sky130_fd_sc_hd__nor2_4 _29883_ (.A(_07539_),
    .B(_07540_),
    .Y(_07547_));
 sky130_vsdinv _29884_ (.A(_07543_),
    .Y(_07548_));
 sky130_fd_sc_hd__o21ai_2 _29885_ (.A1(_07546_),
    .A2(_07547_),
    .B1(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__nand3b_4 _29886_ (.A_N(_07538_),
    .B(_07545_),
    .C(_07549_),
    .Y(_07550_));
 sky130_fd_sc_hd__nand3_4 _29887_ (.A(_07541_),
    .B(_07548_),
    .C(_07544_),
    .Y(_07551_));
 sky130_fd_sc_hd__o21ai_4 _29888_ (.A1(_07546_),
    .A2(_07547_),
    .B1(_07543_),
    .Y(_07552_));
 sky130_fd_sc_hd__nand3_4 _29889_ (.A(_07551_),
    .B(_07538_),
    .C(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__buf_6 _29890_ (.A(\pcpi_mul.rs1[18] ),
    .X(_07554_));
 sky130_fd_sc_hd__nand2_2 _29891_ (.A(_05116_),
    .B(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__buf_6 _29892_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07556_));
 sky130_fd_sc_hd__nand2_2 _29893_ (.A(_05118_),
    .B(_07556_),
    .Y(_07557_));
 sky130_fd_sc_hd__nor2_1 _29894_ (.A(_07555_),
    .B(_07557_),
    .Y(_07558_));
 sky130_fd_sc_hd__and2_1 _29895_ (.A(_07555_),
    .B(_07557_),
    .X(_07559_));
 sky130_vsdinv _29896_ (.A(\pcpi_mul.rs1[17] ),
    .Y(_07560_));
 sky130_fd_sc_hd__buf_2 _29897_ (.A(_07560_),
    .X(_07561_));
 sky130_fd_sc_hd__nor2_4 _29898_ (.A(_05132_),
    .B(net470),
    .Y(_07562_));
 sky130_fd_sc_hd__o21bai_1 _29899_ (.A1(_07558_),
    .A2(_07559_),
    .B1_N(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__or2_1 _29900_ (.A(_07555_),
    .B(_07557_),
    .X(_07564_));
 sky130_fd_sc_hd__nand2_1 _29901_ (.A(_07555_),
    .B(_07557_),
    .Y(_07565_));
 sky130_fd_sc_hd__nand3_2 _29902_ (.A(_07564_),
    .B(_07562_),
    .C(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__nand2_2 _29903_ (.A(_07563_),
    .B(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__nand3_2 _29904_ (.A(_07550_),
    .B(_07553_),
    .C(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__nand2_1 _29905_ (.A(_07550_),
    .B(_07553_),
    .Y(_07569_));
 sky130_vsdinv _29906_ (.A(_07567_),
    .Y(_07570_));
 sky130_fd_sc_hd__nand2_1 _29907_ (.A(_07569_),
    .B(_07570_),
    .Y(_07571_));
 sky130_fd_sc_hd__o2111ai_4 _29908_ (.A1(_07537_),
    .A2(_07352_),
    .B1(_07339_),
    .C1(_07568_),
    .D1(_07571_),
    .Y(_07572_));
 sky130_fd_sc_hd__o21a_1 _29909_ (.A1(_07536_),
    .A2(_07354_),
    .B1(_07572_),
    .X(_07573_));
 sky130_fd_sc_hd__nand3_2 _29910_ (.A(_07570_),
    .B(_07550_),
    .C(_07553_),
    .Y(_07574_));
 sky130_fd_sc_hd__nand2_1 _29911_ (.A(_07569_),
    .B(_07567_),
    .Y(_07575_));
 sky130_fd_sc_hd__o21ai_2 _29912_ (.A1(_07537_),
    .A2(_07352_),
    .B1(_07339_),
    .Y(_07576_));
 sky130_fd_sc_hd__nand3_4 _29913_ (.A(_07574_),
    .B(_07575_),
    .C(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__nor2_1 _29914_ (.A(_07536_),
    .B(_07354_),
    .Y(_07578_));
 sky130_vsdinv _29915_ (.A(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__a21oi_4 _29916_ (.A1(_07572_),
    .A2(_07577_),
    .B1(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__a21oi_4 _29917_ (.A1(_07573_),
    .A2(_07577_),
    .B1(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__o21ai_2 _29918_ (.A1(_07533_),
    .A2(_07535_),
    .B1(_07581_),
    .Y(_07582_));
 sky130_fd_sc_hd__a21o_1 _29919_ (.A1(_07528_),
    .A2(_07531_),
    .B1(_07532_),
    .X(_07583_));
 sky130_fd_sc_hd__nand3_4 _29920_ (.A(_07528_),
    .B(_07532_),
    .C(_07531_),
    .Y(_07584_));
 sky130_fd_sc_hd__a21o_1 _29921_ (.A1(_07572_),
    .A2(_07577_),
    .B1(_07579_),
    .X(_07585_));
 sky130_fd_sc_hd__nand3_1 _29922_ (.A(_07572_),
    .B(_07577_),
    .C(_07579_),
    .Y(_07586_));
 sky130_fd_sc_hd__nand2_1 _29923_ (.A(_07585_),
    .B(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__nand3_2 _29924_ (.A(_07583_),
    .B(_07584_),
    .C(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__nand3_4 _29925_ (.A(_07582_),
    .B(_07254_),
    .C(_07588_),
    .Y(_07589_));
 sky130_vsdinv _29926_ (.A(_07586_),
    .Y(_07590_));
 sky130_fd_sc_hd__o22ai_4 _29927_ (.A1(_07590_),
    .A2(_07580_),
    .B1(_07533_),
    .B2(_07535_),
    .Y(_07591_));
 sky130_vsdinv _29928_ (.A(_07254_),
    .Y(_07592_));
 sky130_fd_sc_hd__nand3_4 _29929_ (.A(_07583_),
    .B(_07584_),
    .C(_07581_),
    .Y(_07593_));
 sky130_fd_sc_hd__nand3_4 _29930_ (.A(_07591_),
    .B(_07592_),
    .C(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__a21bo_2 _29931_ (.A1(_07366_),
    .A2(_07310_),
    .B1_N(_07316_),
    .X(_07595_));
 sky130_fd_sc_hd__a21oi_4 _29932_ (.A1(_07589_),
    .A2(_07594_),
    .B1(_07595_),
    .Y(_07596_));
 sky130_fd_sc_hd__and3_1 _29933_ (.A(_07589_),
    .B(_07594_),
    .C(_07595_),
    .X(_07597_));
 sky130_fd_sc_hd__o22ai_4 _29934_ (.A1(_07498_),
    .A2(_07500_),
    .B1(_07596_),
    .B2(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__nand2_2 _29935_ (.A(_07495_),
    .B(_07496_),
    .Y(_07599_));
 sky130_fd_sc_hd__a21oi_4 _29936_ (.A1(_07599_),
    .A2(_07493_),
    .B1(_07268_),
    .Y(_07600_));
 sky130_fd_sc_hd__a21oi_2 _29937_ (.A1(_07497_),
    .A2(_07600_),
    .B1(_07498_),
    .Y(_07601_));
 sky130_fd_sc_hd__a21o_1 _29938_ (.A1(_07589_),
    .A2(_07594_),
    .B1(_07595_),
    .X(_07602_));
 sky130_fd_sc_hd__nand3_4 _29939_ (.A(_07589_),
    .B(_07594_),
    .C(_07595_),
    .Y(_07603_));
 sky130_fd_sc_hd__nand3_4 _29940_ (.A(_07601_),
    .B(_07602_),
    .C(_07603_),
    .Y(_07604_));
 sky130_vsdinv _29941_ (.A(_07272_),
    .Y(_07605_));
 sky130_fd_sc_hd__nand2_4 _29942_ (.A(_07386_),
    .B(_07605_),
    .Y(_07606_));
 sky130_fd_sc_hd__a21oi_4 _29943_ (.A1(_07598_),
    .A2(_07604_),
    .B1(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__nand2_4 _29944_ (.A(_07600_),
    .B(_07497_),
    .Y(_07608_));
 sky130_fd_sc_hd__nand2_1 _29945_ (.A(_07499_),
    .B(_07271_),
    .Y(_07609_));
 sky130_fd_sc_hd__nand3_4 _29946_ (.A(_07603_),
    .B(_07608_),
    .C(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__o211a_1 _29947_ (.A1(_07596_),
    .A2(_07610_),
    .B1(_07598_),
    .C1(_07606_),
    .X(_07611_));
 sky130_fd_sc_hd__o22ai_4 _29948_ (.A1(_07419_),
    .A2(_07420_),
    .B1(_07607_),
    .B2(_07611_),
    .Y(_07612_));
 sky130_fd_sc_hd__a21o_1 _29949_ (.A1(_07598_),
    .A2(_07604_),
    .B1(_07606_),
    .X(_07613_));
 sky130_fd_sc_hd__nand3_4 _29950_ (.A(_07606_),
    .B(_07598_),
    .C(_07604_),
    .Y(_07614_));
 sky130_fd_sc_hd__nor2_2 _29951_ (.A(_07420_),
    .B(_07419_),
    .Y(_07615_));
 sky130_fd_sc_hd__nand3_4 _29952_ (.A(_07613_),
    .B(_07614_),
    .C(_07615_),
    .Y(_07616_));
 sky130_fd_sc_hd__o21ai_4 _29953_ (.A1(_07396_),
    .A2(_07387_),
    .B1(_07399_),
    .Y(_07617_));
 sky130_fd_sc_hd__a21oi_4 _29954_ (.A1(_07612_),
    .A2(_07616_),
    .B1(_07617_),
    .Y(_07618_));
 sky130_fd_sc_hd__nor2_1 _29955_ (.A(_07396_),
    .B(_07387_),
    .Y(_07619_));
 sky130_fd_sc_hd__o211a_1 _29956_ (.A1(_07388_),
    .A2(_07619_),
    .B1(_07616_),
    .C1(_07612_),
    .X(_07620_));
 sky130_vsdinv _29957_ (.A(_07394_),
    .Y(_07621_));
 sky130_fd_sc_hd__o21ai_2 _29958_ (.A1(_07618_),
    .A2(_07620_),
    .B1(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__a21boi_4 _29959_ (.A1(_07401_),
    .A2(_07409_),
    .B1_N(_07406_),
    .Y(_07623_));
 sky130_fd_sc_hd__a21o_1 _29960_ (.A1(_07612_),
    .A2(_07616_),
    .B1(_07617_),
    .X(_07624_));
 sky130_fd_sc_hd__nand3_4 _29961_ (.A(_07612_),
    .B(_07617_),
    .C(_07616_),
    .Y(_07625_));
 sky130_fd_sc_hd__nand3_2 _29962_ (.A(_07624_),
    .B(_07394_),
    .C(_07625_),
    .Y(_07626_));
 sky130_fd_sc_hd__nand3_4 _29963_ (.A(_07622_),
    .B(_07623_),
    .C(_07626_),
    .Y(_07627_));
 sky130_vsdinv _29964_ (.A(_07389_),
    .Y(_07628_));
 sky130_fd_sc_hd__o22ai_4 _29965_ (.A1(_07392_),
    .A2(_07628_),
    .B1(_07618_),
    .B2(_07620_),
    .Y(_07629_));
 sky130_fd_sc_hd__a21bo_1 _29966_ (.A1(_07409_),
    .A2(_07401_),
    .B1_N(_07406_),
    .X(_07630_));
 sky130_fd_sc_hd__nand3_2 _29967_ (.A(_07624_),
    .B(_07621_),
    .C(_07625_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand3_4 _29968_ (.A(_07629_),
    .B(_07630_),
    .C(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__and2_2 _29969_ (.A(_07627_),
    .B(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__o2111ai_4 _29970_ (.A1(_07188_),
    .A2(_07187_),
    .B1(_07189_),
    .C1(_07414_),
    .D1(_07195_),
    .Y(_07634_));
 sky130_fd_sc_hd__or2_4 _29971_ (.A(_07634_),
    .B(_06585_),
    .X(_07635_));
 sky130_fd_sc_hd__nand3_2 _29972_ (.A(_07184_),
    .B(_07181_),
    .C(_07183_),
    .Y(_07636_));
 sky130_fd_sc_hd__o2bb2ai_2 _29973_ (.A1_N(_07410_),
    .A2_N(_07408_),
    .B1(_07636_),
    .B2(_07413_),
    .Y(_07637_));
 sky130_fd_sc_hd__a31oi_4 _29974_ (.A1(_07195_),
    .A2(_07190_),
    .A3(_07414_),
    .B1(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_4 _29975_ (.A(_07635_),
    .B(_07638_),
    .Y(_07639_));
 sky130_fd_sc_hd__xor2_4 _29976_ (.A(_07633_),
    .B(_07639_),
    .X(_02639_));
 sky130_fd_sc_hd__xor2_4 _29977_ (.A(_07416_),
    .B(_07417_),
    .X(_07640_));
 sky130_fd_sc_hd__o21ai_2 _29978_ (.A1(_07640_),
    .A2(_07607_),
    .B1(_07614_),
    .Y(_07641_));
 sky130_fd_sc_hd__buf_6 _29979_ (.A(_19886_),
    .X(_07642_));
 sky130_fd_sc_hd__a22oi_4 _29980_ (.A1(_05440_),
    .A2(_06283_),
    .B1(_05447_),
    .B2(_07642_),
    .Y(_07643_));
 sky130_fd_sc_hd__nand3_4 _29981_ (.A(_19661_),
    .B(_05588_),
    .C(_06779_),
    .Y(_07644_));
 sky130_fd_sc_hd__nor2_4 _29982_ (.A(_06809_),
    .B(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__nand2_2 _29983_ (.A(_05259_),
    .B(_07322_),
    .Y(_07646_));
 sky130_fd_sc_hd__o21ai_2 _29984_ (.A1(_07643_),
    .A2(_07645_),
    .B1(_07646_),
    .Y(_07647_));
 sky130_fd_sc_hd__o21ai_2 _29985_ (.A1(_07465_),
    .A2(_07461_),
    .B1(_07468_),
    .Y(_07648_));
 sky130_vsdinv _29986_ (.A(_07646_),
    .Y(_07649_));
 sky130_fd_sc_hd__a22o_1 _29987_ (.A1(_06492_),
    .A2(_06283_),
    .B1(_06217_),
    .B2(_07642_),
    .X(_07650_));
 sky130_fd_sc_hd__o211ai_2 _29988_ (.A1(_06810_),
    .A2(_07644_),
    .B1(_07649_),
    .C1(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__nand3_4 _29989_ (.A(_07647_),
    .B(_07648_),
    .C(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__o21ai_2 _29990_ (.A1(_07643_),
    .A2(_07645_),
    .B1(_07649_),
    .Y(_07653_));
 sky130_fd_sc_hd__a21oi_2 _29991_ (.A1(_07466_),
    .A2(_07469_),
    .B1(_07464_),
    .Y(_07654_));
 sky130_fd_sc_hd__o211ai_2 _29992_ (.A1(_06810_),
    .A2(_07644_),
    .B1(_07646_),
    .C1(_07650_),
    .Y(_07655_));
 sky130_fd_sc_hd__nand3_4 _29993_ (.A(_07653_),
    .B(_07654_),
    .C(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__nor2_8 _29994_ (.A(_07508_),
    .B(_07504_),
    .Y(_07657_));
 sky130_fd_sc_hd__o2bb2ai_4 _29995_ (.A1_N(_07652_),
    .A2_N(_07656_),
    .B1(_07501_),
    .B2(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__nor2_2 _29996_ (.A(_07501_),
    .B(_07657_),
    .Y(_07659_));
 sky130_fd_sc_hd__nand3_4 _29997_ (.A(_07656_),
    .B(_07652_),
    .C(_07659_),
    .Y(_07660_));
 sky130_vsdinv _29998_ (.A(_07449_),
    .Y(_07661_));
 sky130_fd_sc_hd__nand2_1 _29999_ (.A(_07453_),
    .B(_07454_),
    .Y(_07662_));
 sky130_fd_sc_hd__o2bb2ai_4 _30000_ (.A1_N(_07460_),
    .A2_N(_07471_),
    .B1(_07661_),
    .B2(_07662_),
    .Y(_07663_));
 sky130_fd_sc_hd__a21oi_4 _30001_ (.A1(_07658_),
    .A2(_07660_),
    .B1(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__nand2_1 _30002_ (.A(_07656_),
    .B(_07659_),
    .Y(_07665_));
 sky130_vsdinv _30003_ (.A(_07652_),
    .Y(_07666_));
 sky130_fd_sc_hd__o211a_1 _30004_ (.A1(_07665_),
    .A2(_07666_),
    .B1(_07658_),
    .C1(_07663_),
    .X(_07667_));
 sky130_fd_sc_hd__and2_2 _30005_ (.A(_07523_),
    .B(_07511_),
    .X(_07668_));
 sky130_fd_sc_hd__o21ai_2 _30006_ (.A1(_07664_),
    .A2(_07667_),
    .B1(_07668_),
    .Y(_07669_));
 sky130_fd_sc_hd__o21ai_2 _30007_ (.A1(_07527_),
    .A2(_07522_),
    .B1(_07530_),
    .Y(_07670_));
 sky130_fd_sc_hd__a21o_1 _30008_ (.A1(_07658_),
    .A2(_07660_),
    .B1(_07663_),
    .X(_07671_));
 sky130_fd_sc_hd__nand3_4 _30009_ (.A(_07663_),
    .B(_07658_),
    .C(_07660_),
    .Y(_07672_));
 sky130_fd_sc_hd__nand3b_4 _30010_ (.A_N(_07668_),
    .B(_07671_),
    .C(_07672_),
    .Y(_07673_));
 sky130_fd_sc_hd__nand3_4 _30011_ (.A(_07669_),
    .B(_07670_),
    .C(_07673_),
    .Y(_07674_));
 sky130_fd_sc_hd__o21bai_2 _30012_ (.A1(_07664_),
    .A2(_07667_),
    .B1_N(_07668_),
    .Y(_07675_));
 sky130_fd_sc_hd__nand2_1 _30013_ (.A(_07530_),
    .B(_07527_),
    .Y(_07676_));
 sky130_fd_sc_hd__nand2_1 _30014_ (.A(_07676_),
    .B(_07529_),
    .Y(_07677_));
 sky130_fd_sc_hd__nand3_2 _30015_ (.A(_07671_),
    .B(_07672_),
    .C(_07668_),
    .Y(_07678_));
 sky130_fd_sc_hd__nand3_4 _30016_ (.A(_07675_),
    .B(_07677_),
    .C(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__nand2_1 _30017_ (.A(_07674_),
    .B(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__a21oi_4 _30018_ (.A1(_07551_),
    .A2(_07552_),
    .B1(_07538_),
    .Y(_07681_));
 sky130_fd_sc_hd__o21ai_2 _30019_ (.A1(_07567_),
    .A2(_07681_),
    .B1(_07553_),
    .Y(_07682_));
 sky130_fd_sc_hd__nand2_4 _30020_ (.A(_05284_),
    .B(_19880_),
    .Y(_07683_));
 sky130_fd_sc_hd__nand2_4 _30021_ (.A(_05201_),
    .B(_07050_),
    .Y(_07684_));
 sky130_fd_sc_hd__or2_2 _30022_ (.A(_07683_),
    .B(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__buf_6 _30023_ (.A(\pcpi_mul.rs1[21] ),
    .X(_07686_));
 sky130_fd_sc_hd__nand2_4 _30024_ (.A(net495),
    .B(_07686_),
    .Y(_07687_));
 sky130_vsdinv _30025_ (.A(_07687_),
    .Y(_07688_));
 sky130_fd_sc_hd__nand2_2 _30026_ (.A(_07683_),
    .B(_07684_),
    .Y(_07689_));
 sky130_fd_sc_hd__nand3_4 _30027_ (.A(_07685_),
    .B(_07688_),
    .C(_07689_),
    .Y(_07690_));
 sky130_fd_sc_hd__a21o_1 _30028_ (.A1(_07548_),
    .A2(_07544_),
    .B1(_07547_),
    .X(_07691_));
 sky130_fd_sc_hd__a22oi_4 _30029_ (.A1(_05197_),
    .A2(_06803_),
    .B1(_05562_),
    .B2(_07343_),
    .Y(_07692_));
 sky130_fd_sc_hd__nor2_8 _30030_ (.A(_07683_),
    .B(_07684_),
    .Y(_07693_));
 sky130_fd_sc_hd__o21ai_2 _30031_ (.A1(_07692_),
    .A2(_07693_),
    .B1(_07687_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand3_4 _30032_ (.A(_07690_),
    .B(_07691_),
    .C(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__nand3_2 _30033_ (.A(_07685_),
    .B(_07687_),
    .C(_07689_),
    .Y(_07696_));
 sky130_fd_sc_hd__a21oi_2 _30034_ (.A1(_07548_),
    .A2(_07544_),
    .B1(_07547_),
    .Y(_07697_));
 sky130_fd_sc_hd__o21ai_2 _30035_ (.A1(_07692_),
    .A2(_07693_),
    .B1(_07688_),
    .Y(_07698_));
 sky130_fd_sc_hd__nand3_4 _30036_ (.A(_07696_),
    .B(_07697_),
    .C(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__nand2_1 _30037_ (.A(_07695_),
    .B(_07699_),
    .Y(_07700_));
 sky130_fd_sc_hd__buf_6 _30038_ (.A(\pcpi_mul.rs1[20] ),
    .X(_07701_));
 sky130_fd_sc_hd__buf_6 _30039_ (.A(\pcpi_mul.rs1[19] ),
    .X(_07702_));
 sky130_fd_sc_hd__nand2_2 _30040_ (.A(_05266_),
    .B(_07702_),
    .Y(_07703_));
 sky130_fd_sc_hd__a21o_1 _30041_ (.A1(_05239_),
    .A2(_07701_),
    .B1(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__buf_6 _30042_ (.A(_07542_),
    .X(_07705_));
 sky130_fd_sc_hd__nand3_4 _30043_ (.A(_07703_),
    .B(_05239_),
    .C(_07705_),
    .Y(_07706_));
 sky130_fd_sc_hd__nand2_2 _30044_ (.A(_05670_),
    .B(_07346_),
    .Y(_07707_));
 sky130_fd_sc_hd__a21o_1 _30045_ (.A1(_07704_),
    .A2(_07706_),
    .B1(_07707_),
    .X(_07708_));
 sky130_fd_sc_hd__nand3_1 _30046_ (.A(_07704_),
    .B(_07707_),
    .C(_07706_),
    .Y(_07709_));
 sky130_fd_sc_hd__nand2_2 _30047_ (.A(_07708_),
    .B(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__nand2_2 _30048_ (.A(_07700_),
    .B(_07710_),
    .Y(_07711_));
 sky130_fd_sc_hd__a21oi_4 _30049_ (.A1(_07704_),
    .A2(_07706_),
    .B1(_07707_),
    .Y(_07712_));
 sky130_fd_sc_hd__and3_2 _30050_ (.A(_07704_),
    .B(_07707_),
    .C(_07706_),
    .X(_07713_));
 sky130_fd_sc_hd__nor2_8 _30051_ (.A(_07712_),
    .B(_07713_),
    .Y(_07714_));
 sky130_fd_sc_hd__nand3_4 _30052_ (.A(_07714_),
    .B(_07695_),
    .C(_07699_),
    .Y(_07715_));
 sky130_fd_sc_hd__nand3_4 _30053_ (.A(_07682_),
    .B(_07711_),
    .C(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__nand2_2 _30054_ (.A(_07566_),
    .B(_07564_),
    .Y(_07717_));
 sky130_vsdinv _30055_ (.A(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__a21oi_1 _30056_ (.A1(_07711_),
    .A2(_07715_),
    .B1(_07682_),
    .Y(_07719_));
 sky130_fd_sc_hd__nor2_1 _30057_ (.A(_07718_),
    .B(_07719_),
    .Y(_07720_));
 sky130_fd_sc_hd__and2_1 _30058_ (.A(_07553_),
    .B(_07567_),
    .X(_07721_));
 sky130_fd_sc_hd__a21oi_2 _30059_ (.A1(_07695_),
    .A2(_07699_),
    .B1(_07714_),
    .Y(_07722_));
 sky130_fd_sc_hd__o21a_1 _30060_ (.A1(_07692_),
    .A2(_07693_),
    .B1(_07687_),
    .X(_07723_));
 sky130_fd_sc_hd__o31ai_1 _30061_ (.A1(_07687_),
    .A2(_07692_),
    .A3(_07693_),
    .B1(_07691_),
    .Y(_07724_));
 sky130_fd_sc_hd__o211a_1 _30062_ (.A1(_07723_),
    .A2(_07724_),
    .B1(_07699_),
    .C1(_07714_),
    .X(_07725_));
 sky130_fd_sc_hd__o22ai_4 _30063_ (.A1(_07681_),
    .A2(_07721_),
    .B1(_07722_),
    .B2(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__a21oi_4 _30064_ (.A1(_07726_),
    .A2(_07716_),
    .B1(_07717_),
    .Y(_07727_));
 sky130_fd_sc_hd__a21oi_2 _30065_ (.A1(_07716_),
    .A2(_07720_),
    .B1(_07727_),
    .Y(_07728_));
 sky130_fd_sc_hd__nand2_1 _30066_ (.A(_07680_),
    .B(_07728_),
    .Y(_07729_));
 sky130_fd_sc_hd__a21o_1 _30067_ (.A1(_07726_),
    .A2(_07716_),
    .B1(_07717_),
    .X(_07730_));
 sky130_fd_sc_hd__nand3_2 _30068_ (.A(_07726_),
    .B(_07716_),
    .C(_07717_),
    .Y(_07731_));
 sky130_fd_sc_hd__nand2_2 _30069_ (.A(_07730_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__nand3_2 _30070_ (.A(_07732_),
    .B(_07674_),
    .C(_07679_),
    .Y(_07733_));
 sky130_fd_sc_hd__nand3_4 _30071_ (.A(_07729_),
    .B(_07496_),
    .C(_07733_),
    .Y(_07734_));
 sky130_vsdinv _30072_ (.A(_07731_),
    .Y(_07735_));
 sky130_fd_sc_hd__o2bb2ai_2 _30073_ (.A1_N(_07679_),
    .A2_N(_07674_),
    .B1(_07727_),
    .B2(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__nand3_2 _30074_ (.A(_07728_),
    .B(_07674_),
    .C(_07679_),
    .Y(_07737_));
 sky130_fd_sc_hd__nand3_4 _30075_ (.A(_07736_),
    .B(_07737_),
    .C(_07480_),
    .Y(_07738_));
 sky130_fd_sc_hd__clkbuf_4 _30076_ (.A(_07738_),
    .X(_07739_));
 sky130_fd_sc_hd__nand2_4 _30077_ (.A(_07593_),
    .B(_07584_),
    .Y(_07740_));
 sky130_fd_sc_hd__a21oi_4 _30078_ (.A1(_07734_),
    .A2(_07739_),
    .B1(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__nand3_4 _30079_ (.A(_07734_),
    .B(_07738_),
    .C(_07740_),
    .Y(_07742_));
 sky130_fd_sc_hd__clkbuf_4 _30080_ (.A(\pcpi_mul.rs2[17] ),
    .X(_07743_));
 sky130_fd_sc_hd__buf_6 _30081_ (.A(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__a22oi_4 _30082_ (.A1(_07744_),
    .A2(_05374_),
    .B1(_06921_),
    .B2(_05383_),
    .Y(_07745_));
 sky130_fd_sc_hd__nand3_4 _30083_ (.A(_07743_),
    .B(_19634_),
    .C(_19916_),
    .Y(_07746_));
 sky130_fd_sc_hd__nor2_4 _30084_ (.A(_07200_),
    .B(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__nand2_2 _30085_ (.A(_19640_),
    .B(_05277_),
    .Y(_07748_));
 sky130_vsdinv _30086_ (.A(_07748_),
    .Y(_07749_));
 sky130_fd_sc_hd__o21ai_2 _30087_ (.A1(_07745_),
    .A2(_07747_),
    .B1(_07749_),
    .Y(_07750_));
 sky130_fd_sc_hd__o21ai_1 _30088_ (.A1(_07483_),
    .A2(_07487_),
    .B1(_07482_),
    .Y(_07751_));
 sky130_fd_sc_hd__nand2_2 _30089_ (.A(_07751_),
    .B(_07488_),
    .Y(_07752_));
 sky130_fd_sc_hd__a22o_2 _30090_ (.A1(_19631_),
    .A2(_05224_),
    .B1(_07428_),
    .B2(_05553_),
    .X(_07753_));
 sky130_fd_sc_hd__o211ai_4 _30091_ (.A1(_07426_),
    .A2(_07746_),
    .B1(_07748_),
    .C1(_07753_),
    .Y(_07754_));
 sky130_fd_sc_hd__nand3_1 _30092_ (.A(_07750_),
    .B(_07752_),
    .C(_07754_),
    .Y(_07755_));
 sky130_fd_sc_hd__o21ai_2 _30093_ (.A1(_07745_),
    .A2(_07747_),
    .B1(_07748_),
    .Y(_07756_));
 sky130_fd_sc_hd__buf_6 _30094_ (.A(_19620_),
    .X(_07757_));
 sky130_fd_sc_hd__clkbuf_8 _30095_ (.A(_07258_),
    .X(_07758_));
 sky130_fd_sc_hd__buf_6 _30096_ (.A(_05105_),
    .X(_07759_));
 sky130_fd_sc_hd__a22oi_4 _30097_ (.A1(_07757_),
    .A2(_05198_),
    .B1(_07758_),
    .B2(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__o21ai_2 _30098_ (.A1(_07482_),
    .A2(_07760_),
    .B1(_07485_),
    .Y(_07761_));
 sky130_fd_sc_hd__o211ai_2 _30099_ (.A1(_07426_),
    .A2(_07746_),
    .B1(_07749_),
    .C1(_07753_),
    .Y(_07762_));
 sky130_fd_sc_hd__nand3_4 _30100_ (.A(_07756_),
    .B(_07761_),
    .C(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__o21ai_2 _30101_ (.A1(_07427_),
    .A2(_07423_),
    .B1(_07429_),
    .Y(_07764_));
 sky130_vsdinv _30102_ (.A(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__a21o_2 _30103_ (.A1(_07755_),
    .A2(_07763_),
    .B1(_07765_),
    .X(_07766_));
 sky130_fd_sc_hd__a31oi_4 _30104_ (.A1(_07750_),
    .A2(_07752_),
    .A3(_07754_),
    .B1(_07764_),
    .Y(_07767_));
 sky130_fd_sc_hd__nand2_4 _30105_ (.A(_07767_),
    .B(_07763_),
    .Y(_07768_));
 sky130_fd_sc_hd__nand2_1 _30106_ (.A(_07434_),
    .B(_07436_),
    .Y(_07769_));
 sky130_fd_sc_hd__nand2_4 _30107_ (.A(_07769_),
    .B(_07431_),
    .Y(_07770_));
 sky130_fd_sc_hd__a21oi_4 _30108_ (.A1(_07766_),
    .A2(_07768_),
    .B1(_07770_),
    .Y(_07771_));
 sky130_fd_sc_hd__and3_1 _30109_ (.A(_07766_),
    .B(_07770_),
    .C(_07768_),
    .X(_07772_));
 sky130_fd_sc_hd__a21oi_4 _30110_ (.A1(_07451_),
    .A2(_07452_),
    .B1(_07447_),
    .Y(_07773_));
 sky130_fd_sc_hd__nand2_2 _30111_ (.A(_06413_),
    .B(_05480_),
    .Y(_07774_));
 sky130_fd_sc_hd__nand3b_4 _30112_ (.A_N(_07774_),
    .B(_06345_),
    .C(_05958_),
    .Y(_07775_));
 sky130_fd_sc_hd__nand2_2 _30113_ (.A(_19646_),
    .B(_05660_),
    .Y(_07776_));
 sky130_fd_sc_hd__nand2_2 _30114_ (.A(_07774_),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__nand2_2 _30115_ (.A(_07223_),
    .B(_05558_),
    .Y(_07778_));
 sky130_vsdinv _30116_ (.A(_07778_),
    .Y(_07779_));
 sky130_fd_sc_hd__nand3_2 _30117_ (.A(_07775_),
    .B(_07777_),
    .C(_07779_),
    .Y(_07780_));
 sky130_fd_sc_hd__a22oi_4 _30118_ (.A1(_06608_),
    .A2(_05545_),
    .B1(_06610_),
    .B2(_05672_),
    .Y(_07781_));
 sky130_fd_sc_hd__nor2_2 _30119_ (.A(_07774_),
    .B(_07776_),
    .Y(_07782_));
 sky130_fd_sc_hd__o21ai_2 _30120_ (.A1(_07781_),
    .A2(_07782_),
    .B1(_07778_),
    .Y(_07783_));
 sky130_fd_sc_hd__nand3b_4 _30121_ (.A_N(_07773_),
    .B(_07780_),
    .C(_07783_),
    .Y(_07784_));
 sky130_fd_sc_hd__o21ai_2 _30122_ (.A1(_07781_),
    .A2(_07782_),
    .B1(_07779_),
    .Y(_07785_));
 sky130_fd_sc_hd__nand3_2 _30123_ (.A(_07775_),
    .B(_07777_),
    .C(_07778_),
    .Y(_07786_));
 sky130_fd_sc_hd__nand3_4 _30124_ (.A(_07785_),
    .B(_07786_),
    .C(_07773_),
    .Y(_07787_));
 sky130_fd_sc_hd__nand2_1 _30125_ (.A(_07784_),
    .B(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__buf_4 _30126_ (.A(_19900_),
    .X(_07789_));
 sky130_fd_sc_hd__a22oi_4 _30127_ (.A1(_06326_),
    .A2(_07789_),
    .B1(_06024_),
    .B2(_06440_),
    .Y(_07790_));
 sky130_fd_sc_hd__and4_2 _30128_ (.A(_19651_),
    .B(_05735_),
    .C(_06648_),
    .D(_06259_),
    .X(_07791_));
 sky130_fd_sc_hd__nand2_2 _30129_ (.A(_19658_),
    .B(_06115_),
    .Y(_07792_));
 sky130_vsdinv _30130_ (.A(_07792_),
    .Y(_07793_));
 sky130_fd_sc_hd__o21ai_2 _30131_ (.A1(_07790_),
    .A2(_07791_),
    .B1(_07793_),
    .Y(_07794_));
 sky130_fd_sc_hd__nand2_1 _30132_ (.A(_06882_),
    .B(_06259_),
    .Y(_07795_));
 sky130_fd_sc_hd__nand3b_4 _30133_ (.A_N(_07795_),
    .B(_06019_),
    .C(_05774_),
    .Y(_07796_));
 sky130_fd_sc_hd__a22o_1 _30134_ (.A1(_06401_),
    .A2(_06448_),
    .B1(_05882_),
    .B2(_06657_),
    .X(_07797_));
 sky130_fd_sc_hd__nand3_2 _30135_ (.A(_07796_),
    .B(_07797_),
    .C(_07792_),
    .Y(_07798_));
 sky130_fd_sc_hd__nand2_4 _30136_ (.A(_07794_),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__nand2_1 _30137_ (.A(_07788_),
    .B(_07799_),
    .Y(_07800_));
 sky130_vsdinv _30138_ (.A(_07799_),
    .Y(_07801_));
 sky130_fd_sc_hd__nand3_1 _30139_ (.A(_07801_),
    .B(_07787_),
    .C(_07784_),
    .Y(_07802_));
 sky130_fd_sc_hd__nand2_2 _30140_ (.A(_07800_),
    .B(_07802_),
    .Y(_07803_));
 sky130_fd_sc_hd__o21ai_2 _30141_ (.A1(_07771_),
    .A2(_07772_),
    .B1(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__a21boi_2 _30142_ (.A1(_07443_),
    .A2(_07476_),
    .B1_N(_07440_),
    .Y(_07805_));
 sky130_fd_sc_hd__a21o_1 _30143_ (.A1(_07766_),
    .A2(_07768_),
    .B1(_07770_),
    .X(_07806_));
 sky130_fd_sc_hd__nand3_4 _30144_ (.A(_07766_),
    .B(_07770_),
    .C(_07768_),
    .Y(_07807_));
 sky130_fd_sc_hd__nand2_1 _30145_ (.A(_07788_),
    .B(_07801_),
    .Y(_07808_));
 sky130_fd_sc_hd__nand3_2 _30146_ (.A(_07784_),
    .B(_07787_),
    .C(_07799_),
    .Y(_07809_));
 sky130_fd_sc_hd__nand2_2 _30147_ (.A(_07808_),
    .B(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__nand3_2 _30148_ (.A(_07806_),
    .B(_07807_),
    .C(_07810_),
    .Y(_07811_));
 sky130_fd_sc_hd__nand3_4 _30149_ (.A(_07804_),
    .B(_07805_),
    .C(_07811_),
    .Y(_07812_));
 sky130_vsdinv _30150_ (.A(_07809_),
    .Y(_07813_));
 sky130_vsdinv _30151_ (.A(_07808_),
    .Y(_07814_));
 sky130_fd_sc_hd__o22ai_4 _30152_ (.A1(_07813_),
    .A2(_07814_),
    .B1(_07771_),
    .B2(_07772_),
    .Y(_07815_));
 sky130_fd_sc_hd__a21o_1 _30153_ (.A1(_07455_),
    .A2(_07460_),
    .B1(_07471_),
    .X(_07816_));
 sky130_fd_sc_hd__nand2_1 _30154_ (.A(_07816_),
    .B(_07472_),
    .Y(_07817_));
 sky130_fd_sc_hd__a21oi_1 _30155_ (.A1(_07437_),
    .A2(_07439_),
    .B1(_07438_),
    .Y(_07818_));
 sky130_fd_sc_hd__o21ai_2 _30156_ (.A1(_07817_),
    .A2(_07818_),
    .B1(_07440_),
    .Y(_07819_));
 sky130_fd_sc_hd__nand3_2 _30157_ (.A(_07806_),
    .B(_07807_),
    .C(_07803_),
    .Y(_07820_));
 sky130_fd_sc_hd__nand3_4 _30158_ (.A(_07815_),
    .B(_07819_),
    .C(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__buf_4 _30159_ (.A(\pcpi_mul.rs2[20] ),
    .X(_07822_));
 sky130_fd_sc_hd__nand2_2 _30160_ (.A(_07822_),
    .B(_05122_),
    .Y(_07823_));
 sky130_fd_sc_hd__clkbuf_4 _30161_ (.A(_19624_),
    .X(_07824_));
 sky130_fd_sc_hd__buf_6 _30162_ (.A(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__nand3b_4 _30163_ (.A_N(_07823_),
    .B(_07825_),
    .C(_05121_),
    .Y(_07826_));
 sky130_fd_sc_hd__buf_4 _30164_ (.A(_19624_),
    .X(_07827_));
 sky130_fd_sc_hd__buf_6 _30165_ (.A(\pcpi_mul.rs1[2] ),
    .X(_07828_));
 sky130_fd_sc_hd__nand2_1 _30166_ (.A(_07827_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__nand2_1 _30167_ (.A(_07823_),
    .B(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__nand2_2 _30168_ (.A(_07481_),
    .B(_05467_),
    .Y(_07831_));
 sky130_fd_sc_hd__a21o_1 _30169_ (.A1(_07826_),
    .A2(_07830_),
    .B1(_07831_),
    .X(_07832_));
 sky130_vsdinv _30170_ (.A(_19617_),
    .Y(_07833_));
 sky130_fd_sc_hd__nor2_4 _30171_ (.A(_07833_),
    .B(net453),
    .Y(_07834_));
 sky130_vsdinv _30172_ (.A(_07834_),
    .Y(_07835_));
 sky130_fd_sc_hd__nand3_1 _30173_ (.A(_07826_),
    .B(_07831_),
    .C(_07830_),
    .Y(_07836_));
 sky130_fd_sc_hd__and3_1 _30174_ (.A(_07832_),
    .B(_07835_),
    .C(_07836_),
    .X(_07837_));
 sky130_fd_sc_hd__and2_1 _30175_ (.A(_07832_),
    .B(_07836_),
    .X(_07838_));
 sky130_fd_sc_hd__nor2_4 _30176_ (.A(_07835_),
    .B(_07838_),
    .Y(_07839_));
 sky130_fd_sc_hd__or2_4 _30177_ (.A(_07837_),
    .B(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__a21boi_2 _30178_ (.A1(_07812_),
    .A2(_07821_),
    .B1_N(_07840_),
    .Y(_07841_));
 sky130_fd_sc_hd__nand2_2 _30179_ (.A(_07812_),
    .B(_07821_),
    .Y(_07842_));
 sky130_fd_sc_hd__nor2_4 _30180_ (.A(_07840_),
    .B(_07842_),
    .Y(_07843_));
 sky130_fd_sc_hd__o22ai_4 _30181_ (.A1(_07493_),
    .A2(_07599_),
    .B1(_07841_),
    .B2(_07843_),
    .Y(_07844_));
 sky130_fd_sc_hd__nand2_2 _30182_ (.A(_07842_),
    .B(_07840_),
    .Y(_07845_));
 sky130_fd_sc_hd__nand3b_4 _30183_ (.A_N(_07840_),
    .B(_07812_),
    .C(_07821_),
    .Y(_07846_));
 sky130_fd_sc_hd__nand3b_4 _30184_ (.A_N(_07497_),
    .B(_07845_),
    .C(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__nand3_4 _30185_ (.A(_07742_),
    .B(_07844_),
    .C(_07847_),
    .Y(_07848_));
 sky130_fd_sc_hd__nand2_2 _30186_ (.A(_07844_),
    .B(_07847_),
    .Y(_07849_));
 sky130_fd_sc_hd__nor2_1 _30187_ (.A(_07587_),
    .B(_07533_),
    .Y(_07850_));
 sky130_fd_sc_hd__o2bb2ai_2 _30188_ (.A1_N(_07739_),
    .A2_N(_07734_),
    .B1(_07535_),
    .B2(_07850_),
    .Y(_07851_));
 sky130_fd_sc_hd__nand3b_4 _30189_ (.A_N(_07740_),
    .B(_07739_),
    .C(_07734_),
    .Y(_07852_));
 sky130_fd_sc_hd__nand3_4 _30190_ (.A(_07849_),
    .B(_07851_),
    .C(_07852_),
    .Y(_07853_));
 sky130_fd_sc_hd__o21ai_4 _30191_ (.A1(_07741_),
    .A2(_07848_),
    .B1(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__nand3_4 _30192_ (.A(_07854_),
    .B(_07608_),
    .C(_07604_),
    .Y(_07855_));
 sky130_fd_sc_hd__o22ai_4 _30193_ (.A1(_07271_),
    .A2(_07499_),
    .B1(_07596_),
    .B2(_07610_),
    .Y(_07856_));
 sky130_fd_sc_hd__a21o_1 _30194_ (.A1(_07851_),
    .A2(_07852_),
    .B1(_07849_),
    .X(_07857_));
 sky130_fd_sc_hd__nand3_4 _30195_ (.A(_07856_),
    .B(_07853_),
    .C(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__nand2_1 _30196_ (.A(_07589_),
    .B(_07595_),
    .Y(_07859_));
 sky130_fd_sc_hd__nand2_2 _30197_ (.A(_07859_),
    .B(_07594_),
    .Y(_07860_));
 sky130_vsdinv _30198_ (.A(_07573_),
    .Y(_07861_));
 sky130_fd_sc_hd__nand2_4 _30199_ (.A(_07861_),
    .B(_07577_),
    .Y(_07862_));
 sky130_fd_sc_hd__nand2_2 _30200_ (.A(_07860_),
    .B(_07862_),
    .Y(_07863_));
 sky130_vsdinv _30201_ (.A(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__and2_1 _30202_ (.A(_07859_),
    .B(_07594_),
    .X(_07865_));
 sky130_vsdinv _30203_ (.A(_07862_),
    .Y(_07866_));
 sky130_fd_sc_hd__nand2_1 _30204_ (.A(_07865_),
    .B(_07866_),
    .Y(_07867_));
 sky130_vsdinv _30205_ (.A(_07867_),
    .Y(_07868_));
 sky130_fd_sc_hd__o2bb2ai_2 _30206_ (.A1_N(_07855_),
    .A2_N(_07858_),
    .B1(_07864_),
    .B2(_07868_),
    .Y(_07869_));
 sky130_fd_sc_hd__xor2_4 _30207_ (.A(_07862_),
    .B(_07860_),
    .X(_07870_));
 sky130_fd_sc_hd__nand3_4 _30208_ (.A(_07858_),
    .B(_07870_),
    .C(_07855_),
    .Y(_07871_));
 sky130_fd_sc_hd__nand3_4 _30209_ (.A(_07641_),
    .B(_07869_),
    .C(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__nand2_2 _30210_ (.A(_07867_),
    .B(_07863_),
    .Y(_07873_));
 sky130_fd_sc_hd__nand3_2 _30211_ (.A(_07858_),
    .B(_07855_),
    .C(_07873_),
    .Y(_07874_));
 sky130_fd_sc_hd__a21o_1 _30212_ (.A1(_07858_),
    .A2(_07855_),
    .B1(_07873_),
    .X(_07875_));
 sky130_fd_sc_hd__o2111ai_4 _30213_ (.A1(_07640_),
    .A2(_07607_),
    .B1(_07614_),
    .C1(_07874_),
    .D1(_07875_),
    .Y(_07876_));
 sky130_fd_sc_hd__o2bb2ai_4 _30214_ (.A1_N(_07872_),
    .A2_N(_07876_),
    .B1(_07416_),
    .B2(_07418_),
    .Y(_07877_));
 sky130_fd_sc_hd__nand3_4 _30215_ (.A(_07876_),
    .B(_07419_),
    .C(_07872_),
    .Y(_07878_));
 sky130_fd_sc_hd__o21ai_4 _30216_ (.A1(_07394_),
    .A2(_07618_),
    .B1(_07625_),
    .Y(_07879_));
 sky130_fd_sc_hd__a21oi_4 _30217_ (.A1(_07877_),
    .A2(_07878_),
    .B1(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__and3_1 _30218_ (.A(_07641_),
    .B(_07869_),
    .C(_07871_),
    .X(_07881_));
 sky130_fd_sc_hd__nand2_1 _30219_ (.A(_07876_),
    .B(_07419_),
    .Y(_07882_));
 sky130_fd_sc_hd__o211a_2 _30220_ (.A1(_07881_),
    .A2(_07882_),
    .B1(_07877_),
    .C1(_07879_),
    .X(_07883_));
 sky130_fd_sc_hd__nor2_8 _30221_ (.A(_07880_),
    .B(_07883_),
    .Y(_07884_));
 sky130_vsdinv _30222_ (.A(_07627_),
    .Y(_07885_));
 sky130_fd_sc_hd__a31o_1 _30223_ (.A1(_07635_),
    .A2(_07632_),
    .A3(_07638_),
    .B1(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__xnor2_4 _30224_ (.A(_07884_),
    .B(_07886_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _30225_ (.A(_07858_),
    .B(_07873_),
    .Y(_07887_));
 sky130_fd_sc_hd__and2_1 _30226_ (.A(_07731_),
    .B(_07716_),
    .X(_07888_));
 sky130_fd_sc_hd__a21o_1 _30227_ (.A1(_07742_),
    .A2(_07739_),
    .B1(_07888_),
    .X(_07889_));
 sky130_vsdinv _30228_ (.A(_07889_),
    .Y(_07890_));
 sky130_fd_sc_hd__nand3_1 _30229_ (.A(_07742_),
    .B(_07739_),
    .C(_07888_),
    .Y(_07891_));
 sky130_vsdinv _30230_ (.A(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__buf_6 _30231_ (.A(_06017_),
    .X(_07893_));
 sky130_fd_sc_hd__a22oi_4 _30232_ (.A1(_07893_),
    .A2(_05774_),
    .B1(_06335_),
    .B2(_05962_),
    .Y(_07894_));
 sky130_fd_sc_hd__nand2_2 _30233_ (.A(_06017_),
    .B(_05976_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand2_1 _30234_ (.A(_19654_),
    .B(_07502_),
    .Y(_07896_));
 sky130_fd_sc_hd__nor2_1 _30235_ (.A(_07895_),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__nand2_2 _30236_ (.A(_06013_),
    .B(_06283_),
    .Y(_07898_));
 sky130_fd_sc_hd__o21bai_1 _30237_ (.A1(_07894_),
    .A2(_07897_),
    .B1_N(_07898_),
    .Y(_07899_));
 sky130_fd_sc_hd__nand3b_4 _30238_ (.A_N(_07895_),
    .B(_06159_),
    .C(_06116_),
    .Y(_07900_));
 sky130_fd_sc_hd__nand2_1 _30239_ (.A(_07895_),
    .B(_07896_),
    .Y(_07901_));
 sky130_fd_sc_hd__nand3_1 _30240_ (.A(_07900_),
    .B(_07901_),
    .C(_07898_),
    .Y(_07902_));
 sky130_fd_sc_hd__nand2_2 _30241_ (.A(_07899_),
    .B(_07902_),
    .Y(_07903_));
 sky130_vsdinv _30242_ (.A(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__a22oi_4 _30243_ (.A1(_06341_),
    .A2(_05958_),
    .B1(_06422_),
    .B2(_06257_),
    .Y(_07905_));
 sky130_fd_sc_hd__nand2_2 _30244_ (.A(_19643_),
    .B(_19906_),
    .Y(_07906_));
 sky130_fd_sc_hd__nand2_2 _30245_ (.A(_06897_),
    .B(_06826_),
    .Y(_07907_));
 sky130_fd_sc_hd__nor2_4 _30246_ (.A(_07906_),
    .B(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__nand2_2 _30247_ (.A(_19649_),
    .B(_06448_),
    .Y(_07909_));
 sky130_vsdinv _30248_ (.A(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__o21ai_4 _30249_ (.A1(_07905_),
    .A2(_07908_),
    .B1(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__nand3b_4 _30250_ (.A_N(_07906_),
    .B(_06898_),
    .C(_06827_),
    .Y(_07912_));
 sky130_fd_sc_hd__nand2_2 _30251_ (.A(_07906_),
    .B(_07907_),
    .Y(_07913_));
 sky130_fd_sc_hd__nand3_4 _30252_ (.A(_07912_),
    .B(_07909_),
    .C(_07913_),
    .Y(_07914_));
 sky130_fd_sc_hd__o21ai_1 _30253_ (.A1(_07774_),
    .A2(_07776_),
    .B1(_07778_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_2 _30254_ (.A(_07915_),
    .B(_07777_),
    .Y(_07916_));
 sky130_fd_sc_hd__a21o_2 _30255_ (.A1(_07911_),
    .A2(_07914_),
    .B1(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__nand3_4 _30256_ (.A(_07911_),
    .B(_07914_),
    .C(_07916_),
    .Y(_07918_));
 sky130_fd_sc_hd__nand2_2 _30257_ (.A(_07917_),
    .B(_07918_),
    .Y(_07919_));
 sky130_fd_sc_hd__nor2_2 _30258_ (.A(_07904_),
    .B(_07919_),
    .Y(_07920_));
 sky130_fd_sc_hd__and2_1 _30259_ (.A(_07919_),
    .B(_07904_),
    .X(_07921_));
 sky130_fd_sc_hd__a22oi_4 _30260_ (.A1(_06986_),
    .A2(_05553_),
    .B1(_19635_),
    .B2(_05486_),
    .Y(_07922_));
 sky130_fd_sc_hd__buf_4 _30261_ (.A(_19630_),
    .X(_07923_));
 sky130_fd_sc_hd__and4_4 _30262_ (.A(_07923_),
    .B(_06988_),
    .C(_19913_),
    .D(_05271_),
    .X(_07924_));
 sky130_fd_sc_hd__nand2_2 _30263_ (.A(_19640_),
    .B(_19909_),
    .Y(_07925_));
 sky130_fd_sc_hd__o21ai_2 _30264_ (.A1(_07922_),
    .A2(_07924_),
    .B1(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__nand2_1 _30265_ (.A(_07923_),
    .B(_05377_),
    .Y(_07927_));
 sky130_fd_sc_hd__buf_4 _30266_ (.A(_06920_),
    .X(_07928_));
 sky130_fd_sc_hd__nand3b_4 _30267_ (.A_N(_07927_),
    .B(_07928_),
    .C(_05656_),
    .Y(_07929_));
 sky130_vsdinv _30268_ (.A(_07925_),
    .Y(_07930_));
 sky130_fd_sc_hd__a22o_4 _30269_ (.A1(_06986_),
    .A2(_05208_),
    .B1(_06988_),
    .B2(_19913_),
    .X(_07931_));
 sky130_fd_sc_hd__nand3_4 _30270_ (.A(_07929_),
    .B(_07930_),
    .C(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__buf_4 _30271_ (.A(\pcpi_mul.rs2[20] ),
    .X(_07933_));
 sky130_fd_sc_hd__buf_6 _30272_ (.A(_07933_),
    .X(_07934_));
 sky130_fd_sc_hd__a22oi_4 _30273_ (.A1(_07934_),
    .A2(_07759_),
    .B1(_07825_),
    .B2(_05121_),
    .Y(_07935_));
 sky130_fd_sc_hd__o21ai_2 _30274_ (.A1(_07831_),
    .A2(_07935_),
    .B1(_07826_),
    .Y(_07936_));
 sky130_fd_sc_hd__nand3_4 _30275_ (.A(_07926_),
    .B(_07932_),
    .C(_07936_),
    .Y(_07937_));
 sky130_fd_sc_hd__o21ai_2 _30276_ (.A1(_07922_),
    .A2(_07924_),
    .B1(_07930_),
    .Y(_07938_));
 sky130_fd_sc_hd__nand3_4 _30277_ (.A(_07929_),
    .B(_07925_),
    .C(_07931_),
    .Y(_07939_));
 sky130_fd_sc_hd__o21ai_1 _30278_ (.A1(_07823_),
    .A2(_07829_),
    .B1(_07831_),
    .Y(_07940_));
 sky130_fd_sc_hd__nand2_2 _30279_ (.A(_07940_),
    .B(_07830_),
    .Y(_07941_));
 sky130_fd_sc_hd__nand3_4 _30280_ (.A(_07938_),
    .B(_07939_),
    .C(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__nand2_1 _30281_ (.A(_07937_),
    .B(_07942_),
    .Y(_07943_));
 sky130_fd_sc_hd__o21ai_4 _30282_ (.A1(_07749_),
    .A2(_07747_),
    .B1(_07753_),
    .Y(_07944_));
 sky130_fd_sc_hd__nand2_4 _30283_ (.A(_07943_),
    .B(_07944_),
    .Y(_07945_));
 sky130_vsdinv _30284_ (.A(_07944_),
    .Y(_07946_));
 sky130_fd_sc_hd__nand3_4 _30285_ (.A(_07937_),
    .B(_07942_),
    .C(_07946_),
    .Y(_07947_));
 sky130_fd_sc_hd__nand2_1 _30286_ (.A(_07765_),
    .B(_07755_),
    .Y(_07948_));
 sky130_fd_sc_hd__nand2_4 _30287_ (.A(_07948_),
    .B(_07763_),
    .Y(_07949_));
 sky130_fd_sc_hd__a21oi_4 _30288_ (.A1(_07945_),
    .A2(_07947_),
    .B1(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__and3_1 _30289_ (.A(_07926_),
    .B(_07932_),
    .C(_07936_),
    .X(_07951_));
 sky130_fd_sc_hd__nand2_1 _30290_ (.A(_07942_),
    .B(_07946_),
    .Y(_07952_));
 sky130_fd_sc_hd__o211a_2 _30291_ (.A1(_07951_),
    .A2(_07952_),
    .B1(_07949_),
    .C1(_07945_),
    .X(_07953_));
 sky130_fd_sc_hd__o22ai_4 _30292_ (.A1(_07920_),
    .A2(_07921_),
    .B1(_07950_),
    .B2(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__o21ai_2 _30293_ (.A1(_07810_),
    .A2(_07771_),
    .B1(_07807_),
    .Y(_07955_));
 sky130_fd_sc_hd__a21o_1 _30294_ (.A1(_07945_),
    .A2(_07947_),
    .B1(_07949_),
    .X(_07956_));
 sky130_fd_sc_hd__nand3_4 _30295_ (.A(_07945_),
    .B(_07949_),
    .C(_07947_),
    .Y(_07957_));
 sky130_fd_sc_hd__nand2_1 _30296_ (.A(_07919_),
    .B(_07903_),
    .Y(_07958_));
 sky130_fd_sc_hd__nand3_1 _30297_ (.A(_07904_),
    .B(_07917_),
    .C(_07918_),
    .Y(_07959_));
 sky130_fd_sc_hd__nand2_1 _30298_ (.A(_07958_),
    .B(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__nand3_2 _30299_ (.A(_07956_),
    .B(_07957_),
    .C(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand3_4 _30300_ (.A(_07954_),
    .B(_07955_),
    .C(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__o21ai_2 _30301_ (.A1(_07950_),
    .A2(_07953_),
    .B1(_07960_),
    .Y(_07963_));
 sky130_fd_sc_hd__nand2_1 _30302_ (.A(_07810_),
    .B(_07807_),
    .Y(_07964_));
 sky130_fd_sc_hd__nand2_1 _30303_ (.A(_07964_),
    .B(_07806_),
    .Y(_07965_));
 sky130_fd_sc_hd__nand2_2 _30304_ (.A(_07918_),
    .B(_07903_),
    .Y(_07966_));
 sky130_vsdinv _30305_ (.A(_07917_),
    .Y(_07967_));
 sky130_fd_sc_hd__nand2_1 _30306_ (.A(_07919_),
    .B(_07904_),
    .Y(_07968_));
 sky130_fd_sc_hd__o21ai_4 _30307_ (.A1(_07966_),
    .A2(_07967_),
    .B1(_07968_),
    .Y(_07969_));
 sky130_fd_sc_hd__nand3_2 _30308_ (.A(_07956_),
    .B(_07957_),
    .C(_07969_),
    .Y(_07970_));
 sky130_fd_sc_hd__nand3_4 _30309_ (.A(_07963_),
    .B(_07965_),
    .C(_07970_),
    .Y(_07971_));
 sky130_fd_sc_hd__nand2_1 _30310_ (.A(_07933_),
    .B(_19926_),
    .Y(_07972_));
 sky130_fd_sc_hd__nand3b_2 _30311_ (.A_N(_07972_),
    .B(_07758_),
    .C(_05838_),
    .Y(_07973_));
 sky130_fd_sc_hd__nand2_1 _30312_ (.A(_07827_),
    .B(_05146_),
    .Y(_07974_));
 sky130_fd_sc_hd__nand2_1 _30313_ (.A(_07972_),
    .B(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__nand2_2 _30314_ (.A(_07481_),
    .B(_05236_),
    .Y(_07976_));
 sky130_fd_sc_hd__and3_1 _30315_ (.A(_07973_),
    .B(_07975_),
    .C(_07976_),
    .X(_07977_));
 sky130_fd_sc_hd__buf_6 _30316_ (.A(_19620_),
    .X(_07978_));
 sky130_fd_sc_hd__a22oi_4 _30317_ (.A1(_07978_),
    .A2(_19927_),
    .B1(_19625_),
    .B2(_05264_),
    .Y(_07979_));
 sky130_fd_sc_hd__nor2_1 _30318_ (.A(_07972_),
    .B(_07974_),
    .Y(_07980_));
 sky130_fd_sc_hd__nor2_1 _30319_ (.A(_07979_),
    .B(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__nor2_2 _30320_ (.A(_07976_),
    .B(_07981_),
    .Y(_07982_));
 sky130_fd_sc_hd__nor2_1 _30321_ (.A(_07977_),
    .B(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__buf_4 _30322_ (.A(_19610_),
    .X(_07984_));
 sky130_fd_sc_hd__nand2_1 _30323_ (.A(_07984_),
    .B(_05204_),
    .Y(_07985_));
 sky130_fd_sc_hd__nand2_1 _30324_ (.A(_19616_),
    .B(_05281_),
    .Y(_07986_));
 sky130_fd_sc_hd__nor2_2 _30325_ (.A(_07985_),
    .B(_07986_),
    .Y(_07987_));
 sky130_vsdinv _30326_ (.A(_07987_),
    .Y(_07988_));
 sky130_fd_sc_hd__nand2_1 _30327_ (.A(_07985_),
    .B(_07986_),
    .Y(_07989_));
 sky130_fd_sc_hd__nand2_2 _30328_ (.A(_07988_),
    .B(_07989_),
    .Y(_07990_));
 sky130_fd_sc_hd__nand2_2 _30329_ (.A(_07983_),
    .B(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__o21bai_4 _30330_ (.A1(_07977_),
    .A2(_07982_),
    .B1_N(_07990_),
    .Y(_07992_));
 sky130_fd_sc_hd__a21oi_4 _30331_ (.A1(_07991_),
    .A2(_07992_),
    .B1(_07839_),
    .Y(_07993_));
 sky130_fd_sc_hd__and3_2 _30332_ (.A(_07839_),
    .B(_07991_),
    .C(_07992_),
    .X(_07994_));
 sky130_fd_sc_hd__o2bb2ai_2 _30333_ (.A1_N(_07962_),
    .A2_N(_07971_),
    .B1(_07993_),
    .B2(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__nor2_2 _30334_ (.A(_07993_),
    .B(_07994_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand3_4 _30335_ (.A(_07971_),
    .B(_07962_),
    .C(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__a21boi_4 _30336_ (.A1(_07995_),
    .A2(_07997_),
    .B1_N(_07846_),
    .Y(_07998_));
 sky130_fd_sc_hd__and3_2 _30337_ (.A(_07843_),
    .B(_07995_),
    .C(_07997_),
    .X(_07999_));
 sky130_fd_sc_hd__a22oi_4 _30338_ (.A1(_05440_),
    .A2(_06464_),
    .B1(_05404_),
    .B2(_06443_),
    .Y(_08000_));
 sky130_vsdinv _30339_ (.A(\pcpi_mul.rs1[15] ),
    .Y(_08001_));
 sky130_fd_sc_hd__nand3_4 _30340_ (.A(_05450_),
    .B(_06216_),
    .C(_19887_),
    .Y(_08002_));
 sky130_fd_sc_hd__nor2_4 _30341_ (.A(_08001_),
    .B(_08002_),
    .Y(_08003_));
 sky130_fd_sc_hd__nand2_2 _30342_ (.A(_05259_),
    .B(_06798_),
    .Y(_08004_));
 sky130_fd_sc_hd__o21ai_2 _30343_ (.A1(_08000_),
    .A2(_08003_),
    .B1(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__o21ai_2 _30344_ (.A1(_07792_),
    .A2(_07790_),
    .B1(_07796_),
    .Y(_08006_));
 sky130_fd_sc_hd__clkbuf_8 _30345_ (.A(_08001_),
    .X(_08007_));
 sky130_vsdinv _30346_ (.A(_08004_),
    .Y(_08008_));
 sky130_fd_sc_hd__a22o_2 _30347_ (.A1(_05440_),
    .A2(_07642_),
    .B1(_05404_),
    .B2(_06634_),
    .X(_08009_));
 sky130_fd_sc_hd__o211ai_4 _30348_ (.A1(_08007_),
    .A2(_08002_),
    .B1(_08008_),
    .C1(_08009_),
    .Y(_08010_));
 sky130_fd_sc_hd__nand3_4 _30349_ (.A(_08005_),
    .B(_08006_),
    .C(_08010_),
    .Y(_08011_));
 sky130_fd_sc_hd__o21ai_2 _30350_ (.A1(_08000_),
    .A2(_08003_),
    .B1(_08008_),
    .Y(_08012_));
 sky130_fd_sc_hd__a21oi_4 _30351_ (.A1(_07797_),
    .A2(_07793_),
    .B1(_07791_),
    .Y(_08013_));
 sky130_fd_sc_hd__o211ai_4 _30352_ (.A1(_08007_),
    .A2(_08002_),
    .B1(_08004_),
    .C1(_08009_),
    .Y(_08014_));
 sky130_fd_sc_hd__nand3_4 _30353_ (.A(_08012_),
    .B(_08013_),
    .C(_08014_),
    .Y(_08015_));
 sky130_fd_sc_hd__nor2_4 _30354_ (.A(_07649_),
    .B(_07645_),
    .Y(_08016_));
 sky130_fd_sc_hd__o2bb2ai_4 _30355_ (.A1_N(_08011_),
    .A2_N(_08015_),
    .B1(_07643_),
    .B2(_08016_),
    .Y(_08017_));
 sky130_fd_sc_hd__nor2_2 _30356_ (.A(_07643_),
    .B(_08016_),
    .Y(_08018_));
 sky130_fd_sc_hd__nand3_4 _30357_ (.A(_08015_),
    .B(_08011_),
    .C(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand2_2 _30358_ (.A(_07787_),
    .B(_07799_),
    .Y(_08020_));
 sky130_fd_sc_hd__nand2_4 _30359_ (.A(_08020_),
    .B(_07784_),
    .Y(_08021_));
 sky130_fd_sc_hd__a21oi_4 _30360_ (.A1(_08017_),
    .A2(_08019_),
    .B1(_08021_),
    .Y(_08022_));
 sky130_vsdinv _30361_ (.A(_08011_),
    .Y(_08023_));
 sky130_fd_sc_hd__nand2_1 _30362_ (.A(_08015_),
    .B(_08018_),
    .Y(_08024_));
 sky130_fd_sc_hd__o211a_2 _30363_ (.A1(_08023_),
    .A2(_08024_),
    .B1(_08017_),
    .C1(_08021_),
    .X(_08025_));
 sky130_fd_sc_hd__nand2_2 _30364_ (.A(_07665_),
    .B(_07652_),
    .Y(_08026_));
 sky130_fd_sc_hd__o21ai_2 _30365_ (.A1(_08022_),
    .A2(_08025_),
    .B1(_08026_),
    .Y(_08027_));
 sky130_fd_sc_hd__nand2_1 _30366_ (.A(_07672_),
    .B(_07668_),
    .Y(_08028_));
 sky130_fd_sc_hd__nand2_2 _30367_ (.A(_08028_),
    .B(_07671_),
    .Y(_08029_));
 sky130_fd_sc_hd__nand2_2 _30368_ (.A(_08017_),
    .B(_08019_),
    .Y(_08030_));
 sky130_fd_sc_hd__and2_1 _30369_ (.A(_08020_),
    .B(_07784_),
    .X(_08031_));
 sky130_fd_sc_hd__nand2_2 _30370_ (.A(_08030_),
    .B(_08031_),
    .Y(_08032_));
 sky130_fd_sc_hd__nand3_4 _30371_ (.A(_08021_),
    .B(_08017_),
    .C(_08019_),
    .Y(_08033_));
 sky130_vsdinv _30372_ (.A(_08026_),
    .Y(_08034_));
 sky130_fd_sc_hd__nand3_2 _30373_ (.A(_08032_),
    .B(_08033_),
    .C(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__nand3_4 _30374_ (.A(_08027_),
    .B(_08029_),
    .C(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__o21ai_2 _30375_ (.A1(_08022_),
    .A2(_08025_),
    .B1(_08034_),
    .Y(_08037_));
 sky130_fd_sc_hd__o21ai_2 _30376_ (.A1(_07668_),
    .A2(_07664_),
    .B1(_07672_),
    .Y(_08038_));
 sky130_fd_sc_hd__nand3_2 _30377_ (.A(_08032_),
    .B(_08033_),
    .C(_08026_),
    .Y(_08039_));
 sky130_fd_sc_hd__nand3_4 _30378_ (.A(_08037_),
    .B(_08038_),
    .C(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__nand2_1 _30379_ (.A(_08036_),
    .B(_08040_),
    .Y(_08041_));
 sky130_vsdinv _30380_ (.A(\pcpi_mul.rs1[22] ),
    .Y(_08042_));
 sky130_fd_sc_hd__buf_4 _30381_ (.A(_08042_),
    .X(_08043_));
 sky130_fd_sc_hd__clkbuf_2 _30382_ (.A(_08043_),
    .X(_08044_));
 sky130_fd_sc_hd__nand3_4 _30383_ (.A(_05211_),
    .B(_05201_),
    .C(_07554_),
    .Y(_08045_));
 sky130_fd_sc_hd__a22o_2 _30384_ (.A1(_05284_),
    .A2(_19877_),
    .B1(_05366_),
    .B2(_07345_),
    .X(_08046_));
 sky130_fd_sc_hd__o21ai_2 _30385_ (.A1(net470),
    .A2(_08045_),
    .B1(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__o21ai_4 _30386_ (.A1(net474),
    .A2(_08044_),
    .B1(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__nor2_4 _30387_ (.A(_07560_),
    .B(_08045_),
    .Y(_08049_));
 sky130_fd_sc_hd__nor2_8 _30388_ (.A(_04838_),
    .B(_08042_),
    .Y(_08050_));
 sky130_fd_sc_hd__nand3b_4 _30389_ (.A_N(_08049_),
    .B(_08046_),
    .C(_08050_),
    .Y(_08051_));
 sky130_fd_sc_hd__a21o_2 _30390_ (.A1(_07688_),
    .A2(_07689_),
    .B1(_07693_),
    .X(_08052_));
 sky130_fd_sc_hd__a21oi_4 _30391_ (.A1(_08048_),
    .A2(_08051_),
    .B1(_08052_),
    .Y(_08053_));
 sky130_fd_sc_hd__nor2_1 _30392_ (.A(_07687_),
    .B(_07692_),
    .Y(_08054_));
 sky130_fd_sc_hd__o211a_1 _30393_ (.A1(_07693_),
    .A2(_08054_),
    .B1(_08051_),
    .C1(_08048_),
    .X(_08055_));
 sky130_fd_sc_hd__buf_4 _30394_ (.A(\pcpi_mul.rs1[21] ),
    .X(_08056_));
 sky130_fd_sc_hd__nand2_1 _30395_ (.A(_05125_),
    .B(_07542_),
    .Y(_08057_));
 sky130_fd_sc_hd__a21o_1 _30396_ (.A1(_05382_),
    .A2(_08056_),
    .B1(_08057_),
    .X(_08058_));
 sky130_fd_sc_hd__nand2_1 _30397_ (.A(_19682_),
    .B(_19865_),
    .Y(_08059_));
 sky130_fd_sc_hd__a21o_1 _30398_ (.A1(_05161_),
    .A2(_19868_),
    .B1(_08059_),
    .X(_08060_));
 sky130_fd_sc_hd__buf_6 _30399_ (.A(\pcpi_mul.rs1[19] ),
    .X(_08061_));
 sky130_fd_sc_hd__buf_6 _30400_ (.A(_08061_),
    .X(_08062_));
 sky130_fd_sc_hd__nand2_2 _30401_ (.A(_05670_),
    .B(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__a21o_2 _30402_ (.A1(_08058_),
    .A2(_08060_),
    .B1(_08063_),
    .X(_08064_));
 sky130_fd_sc_hd__nand3_4 _30403_ (.A(_08058_),
    .B(_08060_),
    .C(_08063_),
    .Y(_08065_));
 sky130_fd_sc_hd__nand2_4 _30404_ (.A(_08064_),
    .B(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__o21ai_2 _30405_ (.A1(_08053_),
    .A2(_08055_),
    .B1(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__and2_1 _30406_ (.A(_08064_),
    .B(_08065_),
    .X(_08068_));
 sky130_fd_sc_hd__a21o_1 _30407_ (.A1(_08048_),
    .A2(_08051_),
    .B1(_08052_),
    .X(_08069_));
 sky130_fd_sc_hd__nand3_4 _30408_ (.A(_08048_),
    .B(_08051_),
    .C(_08052_),
    .Y(_08070_));
 sky130_fd_sc_hd__nand3_2 _30409_ (.A(_08068_),
    .B(_08069_),
    .C(_08070_),
    .Y(_08071_));
 sky130_fd_sc_hd__a21oi_2 _30410_ (.A1(_07690_),
    .A2(_07694_),
    .B1(_07691_),
    .Y(_08072_));
 sky130_fd_sc_hd__o21ai_2 _30411_ (.A1(_07710_),
    .A2(_08072_),
    .B1(_07695_),
    .Y(_08073_));
 sky130_fd_sc_hd__nand3_4 _30412_ (.A(_08067_),
    .B(_08071_),
    .C(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__o21a_2 _30413_ (.A1(_07710_),
    .A2(_08072_),
    .B1(_07695_),
    .X(_08075_));
 sky130_fd_sc_hd__o21ai_4 _30414_ (.A1(_08053_),
    .A2(_08055_),
    .B1(_08068_),
    .Y(_08076_));
 sky130_fd_sc_hd__nand3_4 _30415_ (.A(_08069_),
    .B(_08066_),
    .C(_08070_),
    .Y(_08077_));
 sky130_vsdinv _30416_ (.A(\pcpi_mul.rs1[20] ),
    .Y(_08078_));
 sky130_fd_sc_hd__clkbuf_4 _30417_ (.A(_08078_),
    .X(_08079_));
 sky130_fd_sc_hd__buf_8 _30418_ (.A(_08079_),
    .X(_08080_));
 sky130_fd_sc_hd__o31a_4 _30419_ (.A1(_05153_),
    .A2(_08080_),
    .A3(_07703_),
    .B1(_07708_),
    .X(_08081_));
 sky130_fd_sc_hd__a31oi_4 _30420_ (.A1(_08075_),
    .A2(_08076_),
    .A3(_08077_),
    .B1(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__nand3_4 _30421_ (.A(_08075_),
    .B(_08076_),
    .C(_08077_),
    .Y(_08083_));
 sky130_fd_sc_hd__a21boi_4 _30422_ (.A1(_08083_),
    .A2(_08074_),
    .B1_N(_08081_),
    .Y(_08084_));
 sky130_fd_sc_hd__a21oi_4 _30423_ (.A1(_08074_),
    .A2(_08082_),
    .B1(_08084_),
    .Y(_08085_));
 sky130_fd_sc_hd__nand2_1 _30424_ (.A(_08041_),
    .B(_08085_),
    .Y(_08086_));
 sky130_fd_sc_hd__nand2_1 _30425_ (.A(_08083_),
    .B(_08074_),
    .Y(_08087_));
 sky130_fd_sc_hd__nor2_4 _30426_ (.A(_08081_),
    .B(_08087_),
    .Y(_08088_));
 sky130_fd_sc_hd__o211ai_4 _30427_ (.A1(_08084_),
    .A2(_08088_),
    .B1(_08036_),
    .C1(_08040_),
    .Y(_08089_));
 sky130_fd_sc_hd__nand3_4 _30428_ (.A(_08086_),
    .B(_07821_),
    .C(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__o2bb2ai_2 _30429_ (.A1_N(_08036_),
    .A2_N(_08040_),
    .B1(_08088_),
    .B2(_08084_),
    .Y(_08091_));
 sky130_fd_sc_hd__nand3_2 _30430_ (.A(_08085_),
    .B(_08036_),
    .C(_08040_),
    .Y(_08092_));
 sky130_vsdinv _30431_ (.A(_07821_),
    .Y(_08093_));
 sky130_fd_sc_hd__nand3_4 _30432_ (.A(_08091_),
    .B(_08092_),
    .C(_08093_),
    .Y(_08094_));
 sky130_vsdinv _30433_ (.A(_07679_),
    .Y(_08095_));
 sky130_fd_sc_hd__o21ai_4 _30434_ (.A1(_07732_),
    .A2(_08095_),
    .B1(_07674_),
    .Y(_08096_));
 sky130_fd_sc_hd__a21oi_2 _30435_ (.A1(_08090_),
    .A2(_08094_),
    .B1(_08096_),
    .Y(_08097_));
 sky130_vsdinv _30436_ (.A(_07674_),
    .Y(_08098_));
 sky130_fd_sc_hd__nor2_1 _30437_ (.A(_07732_),
    .B(_08095_),
    .Y(_08099_));
 sky130_fd_sc_hd__o211a_1 _30438_ (.A1(_08098_),
    .A2(_08099_),
    .B1(_08094_),
    .C1(_08090_),
    .X(_08100_));
 sky130_fd_sc_hd__o22ai_4 _30439_ (.A1(_07998_),
    .A2(_07999_),
    .B1(_08097_),
    .B2(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__a21o_2 _30440_ (.A1(_08090_),
    .A2(_08094_),
    .B1(_08096_),
    .X(_08102_));
 sky130_fd_sc_hd__nand2_2 _30441_ (.A(_07971_),
    .B(_07962_),
    .Y(_08103_));
 sky130_vsdinv _30442_ (.A(_07996_),
    .Y(_08104_));
 sky130_fd_sc_hd__a21oi_2 _30443_ (.A1(_08103_),
    .A2(_08104_),
    .B1(_07846_),
    .Y(_08105_));
 sky130_fd_sc_hd__a21oi_4 _30444_ (.A1(_07997_),
    .A2(_08105_),
    .B1(_07998_),
    .Y(_08106_));
 sky130_fd_sc_hd__nand3_4 _30445_ (.A(_08090_),
    .B(_08094_),
    .C(_08096_),
    .Y(_08107_));
 sky130_fd_sc_hd__nand3_4 _30446_ (.A(_08102_),
    .B(_08106_),
    .C(_08107_),
    .Y(_08108_));
 sky130_fd_sc_hd__nand2_1 _30447_ (.A(_07845_),
    .B(_07846_),
    .Y(_08109_));
 sky130_fd_sc_hd__o22ai_4 _30448_ (.A1(_07497_),
    .A2(_08109_),
    .B1(_07741_),
    .B2(_07848_),
    .Y(_08110_));
 sky130_fd_sc_hd__a21oi_4 _30449_ (.A1(_08101_),
    .A2(_08108_),
    .B1(_08110_),
    .Y(_08111_));
 sky130_fd_sc_hd__nand2_1 _30450_ (.A(_08102_),
    .B(_08106_),
    .Y(_08112_));
 sky130_fd_sc_hd__o211a_2 _30451_ (.A1(_08100_),
    .A2(_08112_),
    .B1(_08101_),
    .C1(_08110_),
    .X(_08113_));
 sky130_fd_sc_hd__o22ai_4 _30452_ (.A1(_07890_),
    .A2(_07892_),
    .B1(_08111_),
    .B2(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand2_1 _30453_ (.A(_08101_),
    .B(_08108_),
    .Y(_08115_));
 sky130_fd_sc_hd__o21a_1 _30454_ (.A1(_07741_),
    .A2(_07848_),
    .B1(_07847_),
    .X(_08116_));
 sky130_fd_sc_hd__nand2_2 _30455_ (.A(_08115_),
    .B(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__nand2_1 _30456_ (.A(_07889_),
    .B(_07891_),
    .Y(_08118_));
 sky130_vsdinv _30457_ (.A(_08118_),
    .Y(_08119_));
 sky130_fd_sc_hd__nand3_4 _30458_ (.A(_08110_),
    .B(_08101_),
    .C(_08108_),
    .Y(_08120_));
 sky130_fd_sc_hd__nand3_4 _30459_ (.A(_08117_),
    .B(_08119_),
    .C(_08120_),
    .Y(_08121_));
 sky130_fd_sc_hd__a22oi_4 _30460_ (.A1(_07855_),
    .A2(_07887_),
    .B1(_08114_),
    .B2(_08121_),
    .Y(_08122_));
 sky130_fd_sc_hd__o21a_1 _30461_ (.A1(_07596_),
    .A2(_07610_),
    .B1(_07608_),
    .X(_08123_));
 sky130_fd_sc_hd__nor2_1 _30462_ (.A(_07854_),
    .B(_08123_),
    .Y(_08124_));
 sky130_fd_sc_hd__a21oi_1 _30463_ (.A1(_08123_),
    .A2(_07854_),
    .B1(_07873_),
    .Y(_08125_));
 sky130_fd_sc_hd__o211a_1 _30464_ (.A1(_08124_),
    .A2(_08125_),
    .B1(_08121_),
    .C1(_08114_),
    .X(_08126_));
 sky130_fd_sc_hd__o21ai_2 _30465_ (.A1(_08122_),
    .A2(_08126_),
    .B1(_07864_),
    .Y(_08127_));
 sky130_fd_sc_hd__a21boi_4 _30466_ (.A1(_07876_),
    .A2(_07419_),
    .B1_N(_07872_),
    .Y(_08128_));
 sky130_vsdinv _30467_ (.A(_07857_),
    .Y(_08129_));
 sky130_fd_sc_hd__nand2_1 _30468_ (.A(_07856_),
    .B(_07853_),
    .Y(_08130_));
 sky130_fd_sc_hd__o2bb2ai_2 _30469_ (.A1_N(_07855_),
    .A2_N(_07870_),
    .B1(_08129_),
    .B2(_08130_),
    .Y(_08131_));
 sky130_fd_sc_hd__a21o_1 _30470_ (.A1(_08114_),
    .A2(_08121_),
    .B1(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__nand3_4 _30471_ (.A(_08114_),
    .B(_08131_),
    .C(_08121_),
    .Y(_08133_));
 sky130_fd_sc_hd__nand3_2 _30472_ (.A(_08132_),
    .B(_07863_),
    .C(_08133_),
    .Y(_08134_));
 sky130_fd_sc_hd__nand3_4 _30473_ (.A(_08127_),
    .B(_08128_),
    .C(_08134_),
    .Y(_08135_));
 sky130_fd_sc_hd__o22ai_4 _30474_ (.A1(_07866_),
    .A2(_07865_),
    .B1(_08122_),
    .B2(_08126_),
    .Y(_08136_));
 sky130_vsdinv _30475_ (.A(_07419_),
    .Y(_08137_));
 sky130_fd_sc_hd__a21oi_1 _30476_ (.A1(_07869_),
    .A2(_07871_),
    .B1(_07641_),
    .Y(_08138_));
 sky130_fd_sc_hd__o21ai_2 _30477_ (.A1(_08137_),
    .A2(_08138_),
    .B1(_07872_),
    .Y(_08139_));
 sky130_fd_sc_hd__nand3_2 _30478_ (.A(_08132_),
    .B(_07864_),
    .C(_08133_),
    .Y(_08140_));
 sky130_fd_sc_hd__nand3_4 _30479_ (.A(_08136_),
    .B(_08139_),
    .C(_08140_),
    .Y(_08141_));
 sky130_fd_sc_hd__nand2_1 _30480_ (.A(_08135_),
    .B(_08141_),
    .Y(_08142_));
 sky130_fd_sc_hd__nand3_2 _30481_ (.A(_07879_),
    .B(_07877_),
    .C(_07878_),
    .Y(_08143_));
 sky130_fd_sc_hd__a21oi_4 _30482_ (.A1(_07632_),
    .A2(_08143_),
    .B1(_07880_),
    .Y(_08144_));
 sky130_fd_sc_hd__and3_1 _30483_ (.A(_07639_),
    .B(_07633_),
    .C(_07884_),
    .X(_08145_));
 sky130_fd_sc_hd__or3_2 _30484_ (.A(_08142_),
    .B(_08144_),
    .C(_08145_),
    .X(_08146_));
 sky130_fd_sc_hd__o21ai_1 _30485_ (.A1(_08144_),
    .A2(_08145_),
    .B1(_08142_),
    .Y(_08147_));
 sky130_fd_sc_hd__nand2_1 _30486_ (.A(_08146_),
    .B(_08147_),
    .Y(_02641_));
 sky130_fd_sc_hd__o21ai_1 _30487_ (.A1(_08144_),
    .A2(_08145_),
    .B1(_08135_),
    .Y(_08148_));
 sky130_vsdinv _30488_ (.A(_07999_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand2_2 _30489_ (.A(_08108_),
    .B(_08149_),
    .Y(_08150_));
 sky130_fd_sc_hd__nand2_2 _30490_ (.A(_19616_),
    .B(_05120_),
    .Y(_08151_));
 sky130_fd_sc_hd__buf_4 _30491_ (.A(_19606_),
    .X(_08152_));
 sky130_fd_sc_hd__buf_6 _30492_ (.A(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__buf_4 _30493_ (.A(\pcpi_mul.rs2[22] ),
    .X(_08154_));
 sky130_fd_sc_hd__buf_6 _30494_ (.A(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__a22oi_4 _30495_ (.A1(_08153_),
    .A2(_19933_),
    .B1(_08155_),
    .B2(_07759_),
    .Y(_08156_));
 sky130_fd_sc_hd__nand2_2 _30496_ (.A(_19611_),
    .B(_05122_),
    .Y(_08157_));
 sky130_fd_sc_hd__nand2_2 _30497_ (.A(_08152_),
    .B(_19932_),
    .Y(_08158_));
 sky130_fd_sc_hd__nor2_4 _30498_ (.A(_08157_),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__or3_4 _30499_ (.A(_08151_),
    .B(_08156_),
    .C(_08159_),
    .X(_08160_));
 sky130_fd_sc_hd__or2_1 _30500_ (.A(_08157_),
    .B(_08158_),
    .X(_08161_));
 sky130_fd_sc_hd__nand2_2 _30501_ (.A(_08157_),
    .B(_08158_),
    .Y(_08162_));
 sky130_fd_sc_hd__nand2_1 _30502_ (.A(_08161_),
    .B(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__nand2_1 _30503_ (.A(_08163_),
    .B(_08151_),
    .Y(_08164_));
 sky130_fd_sc_hd__nand3_4 _30504_ (.A(_08160_),
    .B(_08164_),
    .C(_07987_),
    .Y(_08165_));
 sky130_vsdinv _30505_ (.A(_08151_),
    .Y(_08166_));
 sky130_fd_sc_hd__nand2_1 _30506_ (.A(_08163_),
    .B(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__nand3_2 _30507_ (.A(_08161_),
    .B(_08162_),
    .C(_08151_),
    .Y(_08168_));
 sky130_fd_sc_hd__nand3_4 _30508_ (.A(_08167_),
    .B(_07988_),
    .C(_08168_),
    .Y(_08169_));
 sky130_fd_sc_hd__nand2_2 _30509_ (.A(_19627_),
    .B(_19917_),
    .Y(_08170_));
 sky130_vsdinv _30510_ (.A(_08170_),
    .Y(_08171_));
 sky130_fd_sc_hd__buf_4 _30511_ (.A(_07258_),
    .X(_08172_));
 sky130_fd_sc_hd__a22oi_4 _30512_ (.A1(_07978_),
    .A2(_05264_),
    .B1(_08172_),
    .B2(_05374_),
    .Y(_08173_));
 sky130_fd_sc_hd__buf_4 _30513_ (.A(_19624_),
    .X(_08174_));
 sky130_fd_sc_hd__nand3_4 _30514_ (.A(_07486_),
    .B(_08174_),
    .C(_05359_),
    .Y(_08175_));
 sky130_fd_sc_hd__nor2_1 _30515_ (.A(_07200_),
    .B(_08175_),
    .Y(_08176_));
 sky130_fd_sc_hd__or3_4 _30516_ (.A(_08171_),
    .B(_08173_),
    .C(_08176_),
    .X(_08177_));
 sky130_fd_sc_hd__o21ai_2 _30517_ (.A1(_08173_),
    .A2(_08176_),
    .B1(_08171_),
    .Y(_08178_));
 sky130_fd_sc_hd__nand2_4 _30518_ (.A(_08177_),
    .B(_08178_),
    .Y(_08179_));
 sky130_fd_sc_hd__a21oi_4 _30519_ (.A1(_08165_),
    .A2(_08169_),
    .B1(_08179_),
    .Y(_08180_));
 sky130_vsdinv _30520_ (.A(_07992_),
    .Y(_08181_));
 sky130_fd_sc_hd__nand3_4 _30521_ (.A(_08165_),
    .B(_08179_),
    .C(_08169_),
    .Y(_08182_));
 sky130_fd_sc_hd__nand2_2 _30522_ (.A(_08181_),
    .B(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__nor2_8 _30523_ (.A(_08180_),
    .B(_08183_),
    .Y(_08184_));
 sky130_fd_sc_hd__a21o_1 _30524_ (.A1(_08165_),
    .A2(_08169_),
    .B1(_08179_),
    .X(_08185_));
 sky130_fd_sc_hd__nand2_2 _30525_ (.A(_08185_),
    .B(_08182_),
    .Y(_08186_));
 sky130_vsdinv _30526_ (.A(_08186_),
    .Y(_08187_));
 sky130_fd_sc_hd__nor2_4 _30527_ (.A(_08181_),
    .B(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__clkbuf_8 _30528_ (.A(_05663_),
    .X(_08189_));
 sky130_fd_sc_hd__buf_6 _30529_ (.A(_19630_),
    .X(_08190_));
 sky130_fd_sc_hd__a22oi_4 _30530_ (.A1(_08190_),
    .A2(_05291_),
    .B1(_19635_),
    .B2(_05481_),
    .Y(_08191_));
 sky130_fd_sc_hd__buf_6 _30531_ (.A(\pcpi_mul.rs2[16] ),
    .X(_08192_));
 sky130_fd_sc_hd__nand3_4 _30532_ (.A(_07923_),
    .B(_08192_),
    .C(_05483_),
    .Y(_08193_));
 sky130_fd_sc_hd__nor2_8 _30533_ (.A(_06214_),
    .B(_08193_),
    .Y(_08194_));
 sky130_fd_sc_hd__o22ai_4 _30534_ (.A1(net441),
    .A2(_08189_),
    .B1(_08191_),
    .B2(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__o21ai_2 _30535_ (.A1(_07976_),
    .A2(_07979_),
    .B1(_07973_),
    .Y(_08196_));
 sky130_fd_sc_hd__buf_8 _30536_ (.A(_06214_),
    .X(_08197_));
 sky130_fd_sc_hd__buf_6 _30537_ (.A(_05480_),
    .X(_08198_));
 sky130_fd_sc_hd__a22o_2 _30538_ (.A1(_08190_),
    .A2(_05291_),
    .B1(_07928_),
    .B2(_08198_),
    .X(_08199_));
 sky130_fd_sc_hd__nor2_8 _30539_ (.A(_06433_),
    .B(_05663_),
    .Y(_08200_));
 sky130_fd_sc_hd__o211ai_4 _30540_ (.A1(_08197_),
    .A2(_08193_),
    .B1(_08199_),
    .C1(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__nand3_4 _30541_ (.A(_08195_),
    .B(_08196_),
    .C(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__o21ai_2 _30542_ (.A1(_08191_),
    .A2(_08194_),
    .B1(_08200_),
    .Y(_08203_));
 sky130_fd_sc_hd__o21ai_1 _30543_ (.A1(_07972_),
    .A2(_07974_),
    .B1(_07976_),
    .Y(_08204_));
 sky130_fd_sc_hd__nand2_2 _30544_ (.A(_08204_),
    .B(_07975_),
    .Y(_08205_));
 sky130_fd_sc_hd__o221ai_4 _30545_ (.A1(_06433_),
    .A2(net449),
    .B1(_08197_),
    .B2(_08193_),
    .C1(_08199_),
    .Y(_08206_));
 sky130_fd_sc_hd__nand3_4 _30546_ (.A(_08203_),
    .B(_08205_),
    .C(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__nor2_2 _30547_ (.A(_07930_),
    .B(_07924_),
    .Y(_08208_));
 sky130_fd_sc_hd__o2bb2ai_4 _30548_ (.A1_N(_08202_),
    .A2_N(_08207_),
    .B1(_07922_),
    .B2(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__a21oi_4 _30549_ (.A1(_07931_),
    .A2(_07930_),
    .B1(_07924_),
    .Y(_08210_));
 sky130_vsdinv _30550_ (.A(_08210_),
    .Y(_08211_));
 sky130_fd_sc_hd__nand3_4 _30551_ (.A(_08207_),
    .B(_08211_),
    .C(_08202_),
    .Y(_08212_));
 sky130_fd_sc_hd__nand2_2 _30552_ (.A(_07952_),
    .B(_07937_),
    .Y(_08213_));
 sky130_fd_sc_hd__a21oi_4 _30553_ (.A1(_08209_),
    .A2(_08212_),
    .B1(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__a31oi_2 _30554_ (.A1(_07938_),
    .A2(_07939_),
    .A3(_07941_),
    .B1(_07944_),
    .Y(_08215_));
 sky130_fd_sc_hd__o211a_4 _30555_ (.A1(_07951_),
    .A2(_08215_),
    .B1(_08212_),
    .C1(_08209_),
    .X(_08216_));
 sky130_fd_sc_hd__a21oi_4 _30556_ (.A1(_07910_),
    .A2(_07913_),
    .B1(_07908_),
    .Y(_08217_));
 sky130_fd_sc_hd__a22oi_4 _30557_ (.A1(_06414_),
    .A2(_05673_),
    .B1(_06345_),
    .B2(_06441_),
    .Y(_08218_));
 sky130_fd_sc_hd__buf_2 _30558_ (.A(_06413_),
    .X(_08219_));
 sky130_fd_sc_hd__and4_1 _30559_ (.A(_08219_),
    .B(_06906_),
    .C(_06448_),
    .D(_05796_),
    .X(_08220_));
 sky130_fd_sc_hd__nand2_4 _30560_ (.A(_19649_),
    .B(_06118_),
    .Y(_08221_));
 sky130_fd_sc_hd__o21ai_2 _30561_ (.A1(_08218_),
    .A2(_08220_),
    .B1(_08221_),
    .Y(_08222_));
 sky130_fd_sc_hd__nand2_1 _30562_ (.A(_07007_),
    .B(_06826_),
    .Y(_08223_));
 sky130_fd_sc_hd__nand3b_4 _30563_ (.A_N(_08223_),
    .B(_19647_),
    .C(_05804_),
    .Y(_08224_));
 sky130_vsdinv _30564_ (.A(_08221_),
    .Y(_08225_));
 sky130_fd_sc_hd__a22o_1 _30565_ (.A1(_06414_),
    .A2(_05673_),
    .B1(_06610_),
    .B2(_07789_),
    .X(_08226_));
 sky130_fd_sc_hd__nand3_2 _30566_ (.A(_08224_),
    .B(_08225_),
    .C(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__nand3b_4 _30567_ (.A_N(_08217_),
    .B(_08222_),
    .C(_08227_),
    .Y(_08228_));
 sky130_fd_sc_hd__o21ai_2 _30568_ (.A1(_08218_),
    .A2(_08220_),
    .B1(_08225_),
    .Y(_08229_));
 sky130_fd_sc_hd__nand3_2 _30569_ (.A(_08224_),
    .B(_08221_),
    .C(_08226_),
    .Y(_08230_));
 sky130_fd_sc_hd__nand3_4 _30570_ (.A(_08229_),
    .B(_08230_),
    .C(_08217_),
    .Y(_08231_));
 sky130_fd_sc_hd__nand2_2 _30571_ (.A(_08228_),
    .B(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__a22oi_4 _30572_ (.A1(_06326_),
    .A2(_06288_),
    .B1(_05736_),
    .B2(_06283_),
    .Y(_08233_));
 sky130_fd_sc_hd__nand2_1 _30573_ (.A(\pcpi_mul.rs2[11] ),
    .B(_19893_),
    .Y(_08234_));
 sky130_fd_sc_hd__nand2_2 _30574_ (.A(_06158_),
    .B(_19890_),
    .Y(_08235_));
 sky130_fd_sc_hd__nor2_1 _30575_ (.A(_08234_),
    .B(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__nand2_2 _30576_ (.A(_19658_),
    .B(_06267_),
    .Y(_08237_));
 sky130_fd_sc_hd__o21bai_1 _30577_ (.A1(_08233_),
    .A2(_08236_),
    .B1_N(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__nand3b_2 _30578_ (.A_N(_08234_),
    .B(_06335_),
    .C(_07281_),
    .Y(_08239_));
 sky130_fd_sc_hd__nand2_1 _30579_ (.A(_08234_),
    .B(_08235_),
    .Y(_08240_));
 sky130_fd_sc_hd__nand3_1 _30580_ (.A(_08239_),
    .B(_08240_),
    .C(_08237_),
    .Y(_08241_));
 sky130_fd_sc_hd__nand2_2 _30581_ (.A(_08238_),
    .B(_08241_),
    .Y(_08242_));
 sky130_vsdinv _30582_ (.A(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__nand2_1 _30583_ (.A(_08232_),
    .B(_08243_),
    .Y(_08244_));
 sky130_fd_sc_hd__nand3_1 _30584_ (.A(_08228_),
    .B(_08231_),
    .C(_08242_),
    .Y(_08245_));
 sky130_fd_sc_hd__nand2_2 _30585_ (.A(_08244_),
    .B(_08245_),
    .Y(_08246_));
 sky130_fd_sc_hd__o21ai_2 _30586_ (.A1(_08214_),
    .A2(_08216_),
    .B1(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__a21o_1 _30587_ (.A1(_08209_),
    .A2(_08212_),
    .B1(_08213_),
    .X(_08248_));
 sky130_fd_sc_hd__nand3_2 _30588_ (.A(_08213_),
    .B(_08209_),
    .C(_08212_),
    .Y(_08249_));
 sky130_fd_sc_hd__nand2_1 _30589_ (.A(_08232_),
    .B(_08242_),
    .Y(_08250_));
 sky130_fd_sc_hd__nand3_2 _30590_ (.A(_08243_),
    .B(_08228_),
    .C(_08231_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_4 _30591_ (.A(_08250_),
    .B(_08251_),
    .Y(_08252_));
 sky130_fd_sc_hd__nand3_2 _30592_ (.A(_08248_),
    .B(_08249_),
    .C(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__nand3_4 _30593_ (.A(_08247_),
    .B(_07994_),
    .C(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__nor2_2 _30594_ (.A(_08242_),
    .B(_08232_),
    .Y(_08255_));
 sky130_fd_sc_hd__and2_1 _30595_ (.A(_08232_),
    .B(_08242_),
    .X(_08256_));
 sky130_fd_sc_hd__o22ai_4 _30596_ (.A1(_08255_),
    .A2(_08256_),
    .B1(_08214_),
    .B2(_08216_),
    .Y(_08257_));
 sky130_fd_sc_hd__nand2_1 _30597_ (.A(_07991_),
    .B(_07992_),
    .Y(_08258_));
 sky130_fd_sc_hd__or2b_1 _30598_ (.A(_08258_),
    .B_N(_07839_),
    .X(_08259_));
 sky130_fd_sc_hd__nand3_2 _30599_ (.A(_08248_),
    .B(_08249_),
    .C(_08246_),
    .Y(_08260_));
 sky130_fd_sc_hd__nand3_4 _30600_ (.A(_08257_),
    .B(_08259_),
    .C(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__o21ai_4 _30601_ (.A1(_07950_),
    .A2(_07969_),
    .B1(_07957_),
    .Y(_08262_));
 sky130_fd_sc_hd__a21oi_4 _30602_ (.A1(_08254_),
    .A2(_08261_),
    .B1(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__nor2_1 _30603_ (.A(_07950_),
    .B(_07969_),
    .Y(_08264_));
 sky130_fd_sc_hd__o211a_4 _30604_ (.A1(_07953_),
    .A2(_08264_),
    .B1(_08261_),
    .C1(_08254_),
    .X(_08265_));
 sky130_fd_sc_hd__o22ai_4 _30605_ (.A1(_08184_),
    .A2(_08188_),
    .B1(_08263_),
    .B2(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__nand2_2 _30606_ (.A(_08254_),
    .B(_08261_),
    .Y(_08267_));
 sky130_vsdinv _30607_ (.A(_08262_),
    .Y(_08268_));
 sky130_fd_sc_hd__nand2_1 _30608_ (.A(_08267_),
    .B(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__nor2_2 _30609_ (.A(_08184_),
    .B(_08188_),
    .Y(_08270_));
 sky130_fd_sc_hd__nand3_4 _30610_ (.A(_08254_),
    .B(_08261_),
    .C(_08262_),
    .Y(_08271_));
 sky130_fd_sc_hd__nand3_4 _30611_ (.A(_08269_),
    .B(_08270_),
    .C(_08271_),
    .Y(_08272_));
 sky130_vsdinv _30612_ (.A(_07997_),
    .Y(_08273_));
 sky130_fd_sc_hd__a21oi_4 _30613_ (.A1(_08266_),
    .A2(_08272_),
    .B1(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__nor2_4 _30614_ (.A(_07992_),
    .B(_08187_),
    .Y(_08275_));
 sky130_fd_sc_hd__nor2_4 _30615_ (.A(_08181_),
    .B(_08186_),
    .Y(_08276_));
 sky130_fd_sc_hd__o2bb2ai_2 _30616_ (.A1_N(_08268_),
    .A2_N(_08267_),
    .B1(_08275_),
    .B2(_08276_),
    .Y(_08277_));
 sky130_fd_sc_hd__o211a_4 _30617_ (.A1(_08265_),
    .A2(_08277_),
    .B1(_08273_),
    .C1(_08266_),
    .X(_08278_));
 sky130_fd_sc_hd__nand2_2 _30618_ (.A(_08033_),
    .B(_08034_),
    .Y(_08279_));
 sky130_fd_sc_hd__buf_4 _30619_ (.A(_06798_),
    .X(_08280_));
 sky130_fd_sc_hd__a22oi_4 _30620_ (.A1(_05832_),
    .A2(_07059_),
    .B1(_06488_),
    .B2(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__nand3_4 _30621_ (.A(_05450_),
    .B(_06216_),
    .C(net497),
    .Y(_08282_));
 sky130_fd_sc_hd__nor2_4 _30622_ (.A(_08001_),
    .B(_08282_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand2_2 _30623_ (.A(_19667_),
    .B(_06783_),
    .Y(_08284_));
 sky130_fd_sc_hd__o21ai_2 _30624_ (.A1(_08281_),
    .A2(_08283_),
    .B1(_08284_),
    .Y(_08285_));
 sky130_vsdinv _30625_ (.A(_08284_),
    .Y(_08286_));
 sky130_fd_sc_hd__a22o_2 _30626_ (.A1(_19662_),
    .A2(_19884_),
    .B1(_06504_),
    .B2(_06799_),
    .X(_08287_));
 sky130_fd_sc_hd__o211ai_4 _30627_ (.A1(_08007_),
    .A2(_08282_),
    .B1(_08286_),
    .C1(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__o21ai_4 _30628_ (.A1(_07898_),
    .A2(_07894_),
    .B1(_07900_),
    .Y(_08289_));
 sky130_fd_sc_hd__nand3_4 _30629_ (.A(_08285_),
    .B(_08288_),
    .C(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__o21ai_2 _30630_ (.A1(_08281_),
    .A2(_08283_),
    .B1(_08286_),
    .Y(_08291_));
 sky130_fd_sc_hd__o21ai_1 _30631_ (.A1(_07895_),
    .A2(_07896_),
    .B1(_07898_),
    .Y(_08292_));
 sky130_fd_sc_hd__nand2_2 _30632_ (.A(_08292_),
    .B(_07901_),
    .Y(_08293_));
 sky130_fd_sc_hd__o211ai_2 _30633_ (.A1(_08007_),
    .A2(_08282_),
    .B1(_08284_),
    .C1(_08287_),
    .Y(_08294_));
 sky130_fd_sc_hd__nand3_4 _30634_ (.A(_08291_),
    .B(_08293_),
    .C(_08294_),
    .Y(_08295_));
 sky130_fd_sc_hd__nor2_4 _30635_ (.A(_08008_),
    .B(_08003_),
    .Y(_08296_));
 sky130_fd_sc_hd__o2bb2ai_4 _30636_ (.A1_N(_08290_),
    .A2_N(_08295_),
    .B1(_08000_),
    .B2(_08296_),
    .Y(_08297_));
 sky130_fd_sc_hd__nor2_2 _30637_ (.A(_08000_),
    .B(_08296_),
    .Y(_08298_));
 sky130_fd_sc_hd__nand3_4 _30638_ (.A(_08290_),
    .B(_08295_),
    .C(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__nand2_4 _30639_ (.A(_07966_),
    .B(_07917_),
    .Y(_08300_));
 sky130_fd_sc_hd__a21oi_4 _30640_ (.A1(_08297_),
    .A2(_08299_),
    .B1(_08300_),
    .Y(_08301_));
 sky130_fd_sc_hd__and3_1 _30641_ (.A(_08285_),
    .B(_08289_),
    .C(_08288_),
    .X(_08302_));
 sky130_fd_sc_hd__nand2_1 _30642_ (.A(_08295_),
    .B(_08298_),
    .Y(_08303_));
 sky130_fd_sc_hd__o211a_1 _30643_ (.A1(_08302_),
    .A2(_08303_),
    .B1(_08297_),
    .C1(_08300_),
    .X(_08304_));
 sky130_fd_sc_hd__nand2_2 _30644_ (.A(_08024_),
    .B(_08011_),
    .Y(_08305_));
 sky130_vsdinv _30645_ (.A(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__o21ai_4 _30646_ (.A1(_08301_),
    .A2(_08304_),
    .B1(_08306_),
    .Y(_08307_));
 sky130_fd_sc_hd__a21o_2 _30647_ (.A1(_08297_),
    .A2(_08299_),
    .B1(_08300_),
    .X(_08308_));
 sky130_fd_sc_hd__nand3_4 _30648_ (.A(_08300_),
    .B(_08297_),
    .C(_08299_),
    .Y(_08309_));
 sky130_fd_sc_hd__nand3_4 _30649_ (.A(_08308_),
    .B(_08309_),
    .C(_08305_),
    .Y(_08310_));
 sky130_fd_sc_hd__a22oi_4 _30650_ (.A1(_08032_),
    .A2(_08279_),
    .B1(_08307_),
    .B2(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__a21oi_4 _30651_ (.A1(_08030_),
    .A2(_08031_),
    .B1(_08034_),
    .Y(_08312_));
 sky130_fd_sc_hd__o211a_2 _30652_ (.A1(_08025_),
    .A2(_08312_),
    .B1(_08310_),
    .C1(_08307_),
    .X(_08313_));
 sky130_fd_sc_hd__a21o_1 _30653_ (.A1(_08050_),
    .A2(_08046_),
    .B1(_08049_),
    .X(_08314_));
 sky130_fd_sc_hd__nand2_4 _30654_ (.A(_05284_),
    .B(_07345_),
    .Y(_08315_));
 sky130_fd_sc_hd__nand2_4 _30655_ (.A(_05285_),
    .B(_08061_),
    .Y(_08316_));
 sky130_fd_sc_hd__nor2_8 _30656_ (.A(_08315_),
    .B(_08316_),
    .Y(_08317_));
 sky130_fd_sc_hd__and2_1 _30657_ (.A(_08315_),
    .B(_08316_),
    .X(_08318_));
 sky130_fd_sc_hd__nand2_2 _30658_ (.A(_05290_),
    .B(_19858_),
    .Y(_08319_));
 sky130_fd_sc_hd__o21ai_2 _30659_ (.A1(_08317_),
    .A2(_08318_),
    .B1(_08319_),
    .Y(_08320_));
 sky130_fd_sc_hd__or2_2 _30660_ (.A(_08315_),
    .B(_08316_),
    .X(_08321_));
 sky130_vsdinv _30661_ (.A(_08319_),
    .Y(_08322_));
 sky130_fd_sc_hd__nand2_4 _30662_ (.A(_08315_),
    .B(_08316_),
    .Y(_08323_));
 sky130_fd_sc_hd__nand3_4 _30663_ (.A(_08321_),
    .B(_08322_),
    .C(_08323_),
    .Y(_08324_));
 sky130_fd_sc_hd__nand3_4 _30664_ (.A(_08314_),
    .B(_08320_),
    .C(_08324_),
    .Y(_08325_));
 sky130_fd_sc_hd__o21ai_2 _30665_ (.A1(_08317_),
    .A2(_08318_),
    .B1(_08322_),
    .Y(_08326_));
 sky130_fd_sc_hd__nand3_2 _30666_ (.A(_08321_),
    .B(_08319_),
    .C(_08323_),
    .Y(_08327_));
 sky130_fd_sc_hd__a21oi_4 _30667_ (.A1(_08050_),
    .A2(_08046_),
    .B1(_08049_),
    .Y(_08328_));
 sky130_fd_sc_hd__nand3_4 _30668_ (.A(_08326_),
    .B(_08327_),
    .C(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__nand2_1 _30669_ (.A(_08325_),
    .B(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__buf_4 _30670_ (.A(_19861_),
    .X(_08331_));
 sky130_fd_sc_hd__buf_6 _30671_ (.A(_08331_),
    .X(_08332_));
 sky130_fd_sc_hd__buf_6 _30672_ (.A(_07686_),
    .X(_08333_));
 sky130_fd_sc_hd__nand2_1 _30673_ (.A(_06636_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__a21o_1 _30674_ (.A1(_05235_),
    .A2(_08332_),
    .B1(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__buf_6 _30675_ (.A(_19865_),
    .X(_08336_));
 sky130_fd_sc_hd__buf_6 _30676_ (.A(_19861_),
    .X(_08337_));
 sky130_fd_sc_hd__nand2_1 _30677_ (.A(_05163_),
    .B(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__a21o_1 _30678_ (.A1(_06639_),
    .A2(_08336_),
    .B1(_08338_),
    .X(_08339_));
 sky130_fd_sc_hd__nand2_2 _30679_ (.A(_05157_),
    .B(_19869_),
    .Y(_08340_));
 sky130_fd_sc_hd__a21o_1 _30680_ (.A1(_08335_),
    .A2(_08339_),
    .B1(_08340_),
    .X(_08341_));
 sky130_fd_sc_hd__nand3_2 _30681_ (.A(_08335_),
    .B(_08339_),
    .C(_08340_),
    .Y(_08342_));
 sky130_fd_sc_hd__nand2_2 _30682_ (.A(_08341_),
    .B(_08342_),
    .Y(_08343_));
 sky130_fd_sc_hd__nand2_2 _30683_ (.A(_08330_),
    .B(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__a21oi_2 _30684_ (.A1(_08335_),
    .A2(_08339_),
    .B1(_08340_),
    .Y(_08345_));
 sky130_vsdinv _30685_ (.A(_08342_),
    .Y(_08346_));
 sky130_fd_sc_hd__nor2_4 _30686_ (.A(_08345_),
    .B(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__nand3_4 _30687_ (.A(_08347_),
    .B(_08325_),
    .C(_08329_),
    .Y(_08348_));
 sky130_fd_sc_hd__o21ai_4 _30688_ (.A1(_08066_),
    .A2(_08053_),
    .B1(_08070_),
    .Y(_08349_));
 sky130_fd_sc_hd__a21oi_1 _30689_ (.A1(_08344_),
    .A2(_08348_),
    .B1(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__and3_1 _30690_ (.A(_08344_),
    .B(_08349_),
    .C(_08348_),
    .X(_08351_));
 sky130_fd_sc_hd__or2_2 _30691_ (.A(_08057_),
    .B(_08059_),
    .X(_08352_));
 sky130_fd_sc_hd__nand2_2 _30692_ (.A(_08064_),
    .B(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__o21ai_1 _30693_ (.A1(_08350_),
    .A2(_08351_),
    .B1(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__a21o_1 _30694_ (.A1(_08344_),
    .A2(_08348_),
    .B1(_08349_),
    .X(_08355_));
 sky130_vsdinv _30695_ (.A(_08353_),
    .Y(_08356_));
 sky130_fd_sc_hd__nand3_4 _30696_ (.A(_08344_),
    .B(_08349_),
    .C(_08348_),
    .Y(_08357_));
 sky130_fd_sc_hd__nand3_1 _30697_ (.A(_08355_),
    .B(_08356_),
    .C(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__nand2_2 _30698_ (.A(_08354_),
    .B(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__o21ai_2 _30699_ (.A1(_08311_),
    .A2(_08313_),
    .B1(_08359_),
    .Y(_08360_));
 sky130_fd_sc_hd__nand2_1 _30700_ (.A(_08355_),
    .B(_08353_),
    .Y(_08361_));
 sky130_fd_sc_hd__o21ai_1 _30701_ (.A1(_08350_),
    .A2(_08351_),
    .B1(_08356_),
    .Y(_08362_));
 sky130_fd_sc_hd__o21ai_1 _30702_ (.A1(_08351_),
    .A2(_08361_),
    .B1(_08362_),
    .Y(_08363_));
 sky130_vsdinv _30703_ (.A(_08279_),
    .Y(_08364_));
 sky130_fd_sc_hd__o2bb2ai_4 _30704_ (.A1_N(_08310_),
    .A2_N(_08307_),
    .B1(_08022_),
    .B2(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__o211ai_4 _30705_ (.A1(_08025_),
    .A2(_08312_),
    .B1(_08310_),
    .C1(_08307_),
    .Y(_08366_));
 sky130_fd_sc_hd__nand3_2 _30706_ (.A(_08363_),
    .B(_08365_),
    .C(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__nand3_4 _30707_ (.A(_08360_),
    .B(_07962_),
    .C(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__a21oi_2 _30708_ (.A1(_08355_),
    .A2(_08357_),
    .B1(_08353_),
    .Y(_08369_));
 sky130_fd_sc_hd__nor2_2 _30709_ (.A(_08351_),
    .B(_08361_),
    .Y(_08370_));
 sky130_fd_sc_hd__o22ai_4 _30710_ (.A1(_08369_),
    .A2(_08370_),
    .B1(_08311_),
    .B2(_08313_),
    .Y(_08371_));
 sky130_vsdinv _30711_ (.A(_07962_),
    .Y(_08372_));
 sky130_fd_sc_hd__nand3_2 _30712_ (.A(_08359_),
    .B(_08365_),
    .C(_08366_),
    .Y(_08373_));
 sky130_fd_sc_hd__nand3_4 _30713_ (.A(_08371_),
    .B(_08372_),
    .C(_08373_),
    .Y(_08374_));
 sky130_fd_sc_hd__nand2_2 _30714_ (.A(_08085_),
    .B(_08036_),
    .Y(_08375_));
 sky130_fd_sc_hd__nand2_4 _30715_ (.A(_08375_),
    .B(_08040_),
    .Y(_08376_));
 sky130_fd_sc_hd__a21oi_4 _30716_ (.A1(_08368_),
    .A2(_08374_),
    .B1(_08376_),
    .Y(_08377_));
 sky130_vsdinv _30717_ (.A(_08040_),
    .Y(_08378_));
 sky130_vsdinv _30718_ (.A(_08375_),
    .Y(_08379_));
 sky130_fd_sc_hd__o211a_2 _30719_ (.A1(_08378_),
    .A2(_08379_),
    .B1(_08374_),
    .C1(_08368_),
    .X(_08380_));
 sky130_fd_sc_hd__o22ai_4 _30720_ (.A1(_08274_),
    .A2(_08278_),
    .B1(_08377_),
    .B2(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__nor2_4 _30721_ (.A(_08276_),
    .B(_08275_),
    .Y(_08382_));
 sky130_fd_sc_hd__nor3_4 _30722_ (.A(_08382_),
    .B(_08263_),
    .C(_08265_),
    .Y(_08383_));
 sky130_fd_sc_hd__nand2_2 _30723_ (.A(_08266_),
    .B(_08273_),
    .Y(_08384_));
 sky130_fd_sc_hd__nand3_4 _30724_ (.A(_08368_),
    .B(_08374_),
    .C(_08376_),
    .Y(_08385_));
 sky130_fd_sc_hd__o2bb2ai_4 _30725_ (.A1_N(_08266_),
    .A2_N(_08272_),
    .B1(_08104_),
    .B2(_08103_),
    .Y(_08386_));
 sky130_fd_sc_hd__a21o_2 _30726_ (.A1(_08368_),
    .A2(_08374_),
    .B1(_08376_),
    .X(_08387_));
 sky130_fd_sc_hd__o2111ai_4 _30727_ (.A1(_08383_),
    .A2(_08384_),
    .B1(_08385_),
    .C1(_08386_),
    .D1(_08387_),
    .Y(_08388_));
 sky130_fd_sc_hd__nand3_4 _30728_ (.A(_08150_),
    .B(_08381_),
    .C(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__a21oi_2 _30729_ (.A1(_08267_),
    .A2(_08268_),
    .B1(_08382_),
    .Y(_08390_));
 sky130_fd_sc_hd__a21o_1 _30730_ (.A1(_08271_),
    .A2(_08390_),
    .B1(_08384_),
    .X(_08391_));
 sky130_fd_sc_hd__o211ai_4 _30731_ (.A1(_08377_),
    .A2(_08380_),
    .B1(_08386_),
    .C1(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__o211ai_4 _30732_ (.A1(_08274_),
    .A2(_08278_),
    .B1(_08387_),
    .C1(_08385_),
    .Y(_08393_));
 sky130_fd_sc_hd__a31oi_4 _30733_ (.A1(_08102_),
    .A2(_08106_),
    .A3(_08107_),
    .B1(_07999_),
    .Y(_08394_));
 sky130_fd_sc_hd__nand3_4 _30734_ (.A(_08392_),
    .B(_08393_),
    .C(_08394_),
    .Y(_08395_));
 sky130_vsdinv _30735_ (.A(_08082_),
    .Y(_08396_));
 sky130_fd_sc_hd__nand2_1 _30736_ (.A(_08396_),
    .B(_08074_),
    .Y(_08397_));
 sky130_fd_sc_hd__nand2_1 _30737_ (.A(_08090_),
    .B(_08096_),
    .Y(_08398_));
 sky130_fd_sc_hd__nand2_1 _30738_ (.A(_08398_),
    .B(_08094_),
    .Y(_08399_));
 sky130_vsdinv _30739_ (.A(_08399_),
    .Y(_08400_));
 sky130_fd_sc_hd__nor2_1 _30740_ (.A(_08397_),
    .B(_08400_),
    .Y(_08401_));
 sky130_vsdinv _30741_ (.A(_08397_),
    .Y(_08402_));
 sky130_fd_sc_hd__nor2_1 _30742_ (.A(_08402_),
    .B(_08399_),
    .Y(_08403_));
 sky130_fd_sc_hd__o2bb2ai_2 _30743_ (.A1_N(_08389_),
    .A2_N(_08395_),
    .B1(_08401_),
    .B2(_08403_),
    .Y(_08404_));
 sky130_fd_sc_hd__a21oi_4 _30744_ (.A1(_08117_),
    .A2(_08119_),
    .B1(_08113_),
    .Y(_08405_));
 sky130_fd_sc_hd__nand2_2 _30745_ (.A(_08399_),
    .B(_08397_),
    .Y(_08406_));
 sky130_fd_sc_hd__nand3_2 _30746_ (.A(_08398_),
    .B(_08094_),
    .C(_08402_),
    .Y(_08407_));
 sky130_fd_sc_hd__nand2_2 _30747_ (.A(_08406_),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__nand3_2 _30748_ (.A(_08395_),
    .B(_08389_),
    .C(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__nand3_4 _30749_ (.A(_08404_),
    .B(_08405_),
    .C(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__inv_2 _30750_ (.A(_08406_),
    .Y(_08411_));
 sky130_vsdinv _30751_ (.A(_08407_),
    .Y(_08412_));
 sky130_fd_sc_hd__o2bb2ai_2 _30752_ (.A1_N(_08389_),
    .A2_N(_08395_),
    .B1(_08411_),
    .B2(_08412_),
    .Y(_08413_));
 sky130_vsdinv _30753_ (.A(_08408_),
    .Y(_08414_));
 sky130_fd_sc_hd__nand3_2 _30754_ (.A(_08395_),
    .B(_08389_),
    .C(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__o21ai_2 _30755_ (.A1(_08118_),
    .A2(_08111_),
    .B1(_08120_),
    .Y(_08416_));
 sky130_fd_sc_hd__nand3_4 _30756_ (.A(_08413_),
    .B(_08415_),
    .C(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__a21o_1 _30757_ (.A1(_08410_),
    .A2(_08417_),
    .B1(_07889_),
    .X(_08418_));
 sky130_fd_sc_hd__nand2_1 _30758_ (.A(_08133_),
    .B(_07863_),
    .Y(_08419_));
 sky130_fd_sc_hd__nand2_1 _30759_ (.A(_08419_),
    .B(_08132_),
    .Y(_08420_));
 sky130_fd_sc_hd__nand3_2 _30760_ (.A(_08410_),
    .B(_08417_),
    .C(_07889_),
    .Y(_08421_));
 sky130_fd_sc_hd__nand3_4 _30761_ (.A(_08418_),
    .B(_08420_),
    .C(_08421_),
    .Y(_08422_));
 sky130_fd_sc_hd__o21ai_1 _30762_ (.A1(_07863_),
    .A2(_08122_),
    .B1(_08133_),
    .Y(_08423_));
 sky130_fd_sc_hd__and2_1 _30763_ (.A(_07742_),
    .B(_07739_),
    .X(_08424_));
 sky130_fd_sc_hd__o2bb2ai_1 _30764_ (.A1_N(_08417_),
    .A2_N(_08410_),
    .B1(_07888_),
    .B2(_08424_),
    .Y(_08425_));
 sky130_fd_sc_hd__nand3_2 _30765_ (.A(_08410_),
    .B(_08417_),
    .C(_07890_),
    .Y(_08426_));
 sky130_fd_sc_hd__nand3_1 _30766_ (.A(_08423_),
    .B(_08425_),
    .C(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__nand2_1 _30767_ (.A(_08422_),
    .B(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__a21oi_1 _30768_ (.A1(_08148_),
    .A2(_08141_),
    .B1(_08428_),
    .Y(_08429_));
 sky130_fd_sc_hd__and3_1 _30769_ (.A(_08148_),
    .B(_08141_),
    .C(_08428_),
    .X(_08430_));
 sky130_fd_sc_hd__nor2_1 _30770_ (.A(_08429_),
    .B(_08430_),
    .Y(_02642_));
 sky130_vsdinv _30771_ (.A(_07878_),
    .Y(_08431_));
 sky130_fd_sc_hd__nand2_1 _30772_ (.A(_07879_),
    .B(_07877_),
    .Y(_08432_));
 sky130_fd_sc_hd__a21o_1 _30773_ (.A1(_07877_),
    .A2(_07878_),
    .B1(_07879_),
    .X(_08433_));
 sky130_fd_sc_hd__o2111ai_4 _30774_ (.A1(_08431_),
    .A2(_08432_),
    .B1(_07627_),
    .C1(_07632_),
    .D1(_08433_),
    .Y(_08434_));
 sky130_vsdinv _30775_ (.A(_08426_),
    .Y(_08435_));
 sky130_fd_sc_hd__nand2_1 _30776_ (.A(_08423_),
    .B(_08425_),
    .Y(_08436_));
 sky130_fd_sc_hd__o2111ai_4 _30777_ (.A1(_08435_),
    .A2(_08436_),
    .B1(_08135_),
    .C1(_08141_),
    .D1(_08422_),
    .Y(_08437_));
 sky130_fd_sc_hd__nor3_4 _30778_ (.A(_08434_),
    .B(_08437_),
    .C(_07634_),
    .Y(_08438_));
 sky130_fd_sc_hd__nand2_8 _30779_ (.A(_06584_),
    .B(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__a31oi_4 _30780_ (.A1(_08387_),
    .A2(_08386_),
    .A3(_08385_),
    .B1(_08278_),
    .Y(_08440_));
 sky130_fd_sc_hd__nand2_2 _30781_ (.A(_08306_),
    .B(_08309_),
    .Y(_08441_));
 sky130_fd_sc_hd__a22oi_4 _30782_ (.A1(_19662_),
    .A2(_06799_),
    .B1(_06504_),
    .B2(_07056_),
    .Y(_08442_));
 sky130_fd_sc_hd__nor2_4 _30783_ (.A(net470),
    .B(_08282_),
    .Y(_08443_));
 sky130_fd_sc_hd__nand2_2 _30784_ (.A(_05443_),
    .B(_07345_),
    .Y(_08444_));
 sky130_fd_sc_hd__o21ai_2 _30785_ (.A1(_08442_),
    .A2(_08443_),
    .B1(_08444_),
    .Y(_08445_));
 sky130_fd_sc_hd__o21ai_2 _30786_ (.A1(_08237_),
    .A2(_08233_),
    .B1(_08239_),
    .Y(_08446_));
 sky130_fd_sc_hd__buf_8 _30787_ (.A(_07560_),
    .X(_08447_));
 sky130_vsdinv _30788_ (.A(_08444_),
    .Y(_08448_));
 sky130_fd_sc_hd__a22o_1 _30789_ (.A1(_05832_),
    .A2(_08280_),
    .B1(_05833_),
    .B2(_07343_),
    .X(_08449_));
 sky130_fd_sc_hd__o211ai_2 _30790_ (.A1(_08447_),
    .A2(_08282_),
    .B1(_08448_),
    .C1(_08449_),
    .Y(_08450_));
 sky130_fd_sc_hd__nand3_4 _30791_ (.A(_08445_),
    .B(_08446_),
    .C(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__o21ai_2 _30792_ (.A1(_08442_),
    .A2(_08443_),
    .B1(_08448_),
    .Y(_08452_));
 sky130_fd_sc_hd__o21ai_1 _30793_ (.A1(_08234_),
    .A2(_08235_),
    .B1(_08237_),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_2 _30794_ (.A(_08453_),
    .B(_08240_),
    .Y(_08454_));
 sky130_fd_sc_hd__o211ai_2 _30795_ (.A1(_08447_),
    .A2(_08282_),
    .B1(_08444_),
    .C1(_08449_),
    .Y(_08455_));
 sky130_fd_sc_hd__nand3_4 _30796_ (.A(_08452_),
    .B(_08454_),
    .C(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__nor2_4 _30797_ (.A(_08286_),
    .B(_08283_),
    .Y(_08457_));
 sky130_fd_sc_hd__o2bb2ai_4 _30798_ (.A1_N(_08451_),
    .A2_N(_08456_),
    .B1(_08281_),
    .B2(_08457_),
    .Y(_08458_));
 sky130_fd_sc_hd__nor2_2 _30799_ (.A(_08281_),
    .B(_08457_),
    .Y(_08459_));
 sky130_fd_sc_hd__nand3_4 _30800_ (.A(_08451_),
    .B(_08456_),
    .C(_08459_),
    .Y(_08460_));
 sky130_fd_sc_hd__nand2_1 _30801_ (.A(_08231_),
    .B(_08242_),
    .Y(_08461_));
 sky130_fd_sc_hd__nand2_4 _30802_ (.A(_08461_),
    .B(_08228_),
    .Y(_08462_));
 sky130_fd_sc_hd__a21oi_4 _30803_ (.A1(_08458_),
    .A2(_08460_),
    .B1(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__nand2_1 _30804_ (.A(_08456_),
    .B(_08459_),
    .Y(_08464_));
 sky130_vsdinv _30805_ (.A(_08451_),
    .Y(_08465_));
 sky130_fd_sc_hd__o211a_1 _30806_ (.A1(_08464_),
    .A2(_08465_),
    .B1(_08458_),
    .C1(_08462_),
    .X(_08466_));
 sky130_fd_sc_hd__and2_2 _30807_ (.A(_08303_),
    .B(_08290_),
    .X(_08467_));
 sky130_fd_sc_hd__o21ai_4 _30808_ (.A1(_08463_),
    .A2(_08466_),
    .B1(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__a21o_1 _30809_ (.A1(_08458_),
    .A2(_08460_),
    .B1(_08462_),
    .X(_08469_));
 sky130_fd_sc_hd__nand3_4 _30810_ (.A(_08462_),
    .B(_08458_),
    .C(_08460_),
    .Y(_08470_));
 sky130_fd_sc_hd__nand3b_4 _30811_ (.A_N(_08467_),
    .B(_08469_),
    .C(_08470_),
    .Y(_08471_));
 sky130_fd_sc_hd__a22oi_4 _30812_ (.A1(_08308_),
    .A2(_08441_),
    .B1(_08468_),
    .B2(_08471_),
    .Y(_08472_));
 sky130_fd_sc_hd__nor2_1 _30813_ (.A(_08306_),
    .B(_08301_),
    .Y(_08473_));
 sky130_fd_sc_hd__o211a_2 _30814_ (.A1(_08304_),
    .A2(_08473_),
    .B1(_08471_),
    .C1(_08468_),
    .X(_08474_));
 sky130_fd_sc_hd__nand2_1 _30815_ (.A(_05266_),
    .B(_08331_),
    .Y(_08475_));
 sky130_fd_sc_hd__a21o_1 _30816_ (.A1(_05119_),
    .A2(_19858_),
    .B1(_08475_),
    .X(_08476_));
 sky130_fd_sc_hd__buf_4 _30817_ (.A(\pcpi_mul.rs1[23] ),
    .X(_08477_));
 sky130_fd_sc_hd__nand2_1 _30818_ (.A(_05152_),
    .B(_08477_),
    .Y(_08478_));
 sky130_fd_sc_hd__a21o_1 _30819_ (.A1(_19679_),
    .A2(_08337_),
    .B1(_08478_),
    .X(_08479_));
 sky130_fd_sc_hd__nand2_2 _30820_ (.A(_05670_),
    .B(_08336_),
    .Y(_08480_));
 sky130_fd_sc_hd__nand3_1 _30821_ (.A(_08476_),
    .B(_08479_),
    .C(_08480_),
    .Y(_08481_));
 sky130_vsdinv _30822_ (.A(_08481_),
    .Y(_08482_));
 sky130_fd_sc_hd__a21oi_4 _30823_ (.A1(_08476_),
    .A2(_08479_),
    .B1(_08480_),
    .Y(_08483_));
 sky130_fd_sc_hd__and4_2 _30824_ (.A(_05294_),
    .B(_19672_),
    .C(\pcpi_mul.rs1[20] ),
    .D(_07556_),
    .X(_08484_));
 sky130_fd_sc_hd__buf_4 _30825_ (.A(\pcpi_mul.rs1[20] ),
    .X(_08485_));
 sky130_fd_sc_hd__a22o_2 _30826_ (.A1(_19670_),
    .A2(_07702_),
    .B1(_05358_),
    .B2(_08485_),
    .X(_08486_));
 sky130_vsdinv _30827_ (.A(\pcpi_mul.rs1[24] ),
    .Y(_08487_));
 sky130_fd_sc_hd__nor2_8 _30828_ (.A(_04838_),
    .B(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__nand3b_4 _30829_ (.A_N(_08484_),
    .B(_08486_),
    .C(_08488_),
    .Y(_08489_));
 sky130_fd_sc_hd__a22oi_4 _30830_ (.A1(_05197_),
    .A2(_07325_),
    .B1(_19673_),
    .B2(_19868_),
    .Y(_08490_));
 sky130_fd_sc_hd__o21bai_4 _30831_ (.A1(_08490_),
    .A2(_08484_),
    .B1_N(_08488_),
    .Y(_08491_));
 sky130_fd_sc_hd__a21o_1 _30832_ (.A1(_08322_),
    .A2(_08323_),
    .B1(_08317_),
    .X(_08492_));
 sky130_fd_sc_hd__a21oi_4 _30833_ (.A1(_08489_),
    .A2(_08491_),
    .B1(_08492_),
    .Y(_08493_));
 sky130_fd_sc_hd__a21oi_4 _30834_ (.A1(_08322_),
    .A2(_08323_),
    .B1(_08317_),
    .Y(_08494_));
 sky130_fd_sc_hd__nand2_4 _30835_ (.A(_08489_),
    .B(_08491_),
    .Y(_08495_));
 sky130_fd_sc_hd__nor2_4 _30836_ (.A(_08494_),
    .B(_08495_),
    .Y(_08496_));
 sky130_fd_sc_hd__o22ai_4 _30837_ (.A1(_08482_),
    .A2(_08483_),
    .B1(_08493_),
    .B2(_08496_),
    .Y(_08497_));
 sky130_fd_sc_hd__a21oi_1 _30838_ (.A1(_08320_),
    .A2(_08324_),
    .B1(_08314_),
    .Y(_08498_));
 sky130_fd_sc_hd__o21ai_2 _30839_ (.A1(_08343_),
    .A2(_08498_),
    .B1(_08325_),
    .Y(_08499_));
 sky130_fd_sc_hd__nor2_8 _30840_ (.A(_08483_),
    .B(_08482_),
    .Y(_08500_));
 sky130_fd_sc_hd__nand2_4 _30841_ (.A(_08495_),
    .B(_08494_),
    .Y(_08501_));
 sky130_fd_sc_hd__nand3_4 _30842_ (.A(_08489_),
    .B(_08491_),
    .C(_08492_),
    .Y(_08502_));
 sky130_fd_sc_hd__nand3_4 _30843_ (.A(_08500_),
    .B(_08501_),
    .C(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__nand3_4 _30844_ (.A(_08497_),
    .B(_08499_),
    .C(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__o21ai_4 _30845_ (.A1(_08493_),
    .A2(_08496_),
    .B1(_08500_),
    .Y(_08505_));
 sky130_fd_sc_hd__a21boi_4 _30846_ (.A1(_08347_),
    .A2(_08329_),
    .B1_N(_08325_),
    .Y(_08506_));
 sky130_fd_sc_hd__o211ai_4 _30847_ (.A1(_08482_),
    .A2(_08483_),
    .B1(_08502_),
    .C1(_08501_),
    .Y(_08507_));
 sky130_fd_sc_hd__o21a_2 _30848_ (.A1(_08334_),
    .A2(_08338_),
    .B1(_08341_),
    .X(_08508_));
 sky130_fd_sc_hd__a31oi_4 _30849_ (.A1(_08505_),
    .A2(_08506_),
    .A3(_08507_),
    .B1(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__nand3_4 _30850_ (.A(_08505_),
    .B(_08506_),
    .C(_08507_),
    .Y(_08510_));
 sky130_fd_sc_hd__a21boi_4 _30851_ (.A1(_08510_),
    .A2(_08504_),
    .B1_N(_08508_),
    .Y(_08511_));
 sky130_fd_sc_hd__a21oi_4 _30852_ (.A1(_08504_),
    .A2(_08509_),
    .B1(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__o21ai_2 _30853_ (.A1(_08472_),
    .A2(_08474_),
    .B1(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__a21boi_4 _30854_ (.A1(_08261_),
    .A2(_08262_),
    .B1_N(_08254_),
    .Y(_08514_));
 sky130_fd_sc_hd__nand2_1 _30855_ (.A(_08468_),
    .B(_08471_),
    .Y(_08515_));
 sky130_fd_sc_hd__nand2_1 _30856_ (.A(_08441_),
    .B(_08308_),
    .Y(_08516_));
 sky130_fd_sc_hd__nand2_2 _30857_ (.A(_08515_),
    .B(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__nand3b_4 _30858_ (.A_N(_08516_),
    .B(_08471_),
    .C(_08468_),
    .Y(_08518_));
 sky130_fd_sc_hd__nand2_1 _30859_ (.A(_08510_),
    .B(_08504_),
    .Y(_08519_));
 sky130_fd_sc_hd__nand2_1 _30860_ (.A(_08519_),
    .B(_08508_),
    .Y(_08520_));
 sky130_fd_sc_hd__nand2_1 _30861_ (.A(_08509_),
    .B(_08504_),
    .Y(_08521_));
 sky130_fd_sc_hd__nand2_2 _30862_ (.A(_08520_),
    .B(_08521_),
    .Y(_08522_));
 sky130_fd_sc_hd__nand3_2 _30863_ (.A(_08517_),
    .B(_08518_),
    .C(_08522_),
    .Y(_08523_));
 sky130_fd_sc_hd__nand3_4 _30864_ (.A(_08513_),
    .B(_08514_),
    .C(_08523_),
    .Y(_08524_));
 sky130_fd_sc_hd__nor2_2 _30865_ (.A(_08508_),
    .B(_08519_),
    .Y(_08525_));
 sky130_fd_sc_hd__o22ai_4 _30866_ (.A1(_08525_),
    .A2(_08511_),
    .B1(_08472_),
    .B2(_08474_),
    .Y(_08526_));
 sky130_fd_sc_hd__nand2_1 _30867_ (.A(_08261_),
    .B(_08262_),
    .Y(_08527_));
 sky130_fd_sc_hd__nand2_2 _30868_ (.A(_08527_),
    .B(_08254_),
    .Y(_08528_));
 sky130_fd_sc_hd__nand3_2 _30869_ (.A(_08517_),
    .B(_08512_),
    .C(_08518_),
    .Y(_08529_));
 sky130_fd_sc_hd__nand3_4 _30870_ (.A(_08526_),
    .B(_08528_),
    .C(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__a21oi_4 _30871_ (.A1(_08359_),
    .A2(_08365_),
    .B1(_08313_),
    .Y(_08531_));
 sky130_vsdinv _30872_ (.A(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__a21oi_4 _30873_ (.A1(_08524_),
    .A2(_08530_),
    .B1(_08532_),
    .Y(_08533_));
 sky130_fd_sc_hd__nand2_2 _30874_ (.A(_08524_),
    .B(_08530_),
    .Y(_08534_));
 sky130_fd_sc_hd__nor2_4 _30875_ (.A(_08531_),
    .B(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__nand2_1 _30876_ (.A(_08179_),
    .B(_08169_),
    .Y(_08536_));
 sky130_fd_sc_hd__nand2_1 _30877_ (.A(_08536_),
    .B(_08165_),
    .Y(_08537_));
 sky130_fd_sc_hd__nor2_2 _30878_ (.A(_08151_),
    .B(_08156_),
    .Y(_08538_));
 sky130_fd_sc_hd__buf_4 _30879_ (.A(\pcpi_mul.rs2[23] ),
    .X(_08539_));
 sky130_fd_sc_hd__nand2_2 _30880_ (.A(_08539_),
    .B(_05105_),
    .Y(_08540_));
 sky130_fd_sc_hd__buf_8 _30881_ (.A(_19611_),
    .X(_08541_));
 sky130_fd_sc_hd__nand3b_4 _30882_ (.A_N(_08540_),
    .B(_08541_),
    .C(_05230_),
    .Y(_08542_));
 sky130_fd_sc_hd__nand2_2 _30883_ (.A(_07984_),
    .B(_05127_),
    .Y(_08543_));
 sky130_fd_sc_hd__nand2_2 _30884_ (.A(_08540_),
    .B(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__buf_4 _30885_ (.A(\pcpi_mul.rs2[21] ),
    .X(_08545_));
 sky130_fd_sc_hd__nand2_2 _30886_ (.A(_08545_),
    .B(_05467_),
    .Y(_08546_));
 sky130_vsdinv _30887_ (.A(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand3_2 _30888_ (.A(_08542_),
    .B(_08544_),
    .C(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__buf_4 _30889_ (.A(_19606_),
    .X(_08549_));
 sky130_fd_sc_hd__buf_6 _30890_ (.A(_08154_),
    .X(_08550_));
 sky130_fd_sc_hd__a22oi_4 _30891_ (.A1(_08549_),
    .A2(_05199_),
    .B1(_08550_),
    .B2(_05230_),
    .Y(_08551_));
 sky130_fd_sc_hd__nor2_4 _30892_ (.A(_08540_),
    .B(_08543_),
    .Y(_08552_));
 sky130_fd_sc_hd__o21ai_2 _30893_ (.A1(_08551_),
    .A2(_08552_),
    .B1(_08546_),
    .Y(_08553_));
 sky130_fd_sc_hd__o211ai_4 _30894_ (.A1(_08159_),
    .A2(_08538_),
    .B1(_08548_),
    .C1(_08553_),
    .Y(_08554_));
 sky130_fd_sc_hd__o21ai_2 _30895_ (.A1(_08551_),
    .A2(_08552_),
    .B1(_08547_),
    .Y(_08555_));
 sky130_fd_sc_hd__nand3_2 _30896_ (.A(_08542_),
    .B(_08544_),
    .C(_08546_),
    .Y(_08556_));
 sky130_fd_sc_hd__a21oi_2 _30897_ (.A1(_08166_),
    .A2(_08162_),
    .B1(_08159_),
    .Y(_08557_));
 sky130_fd_sc_hd__nand3_4 _30898_ (.A(_08555_),
    .B(_08556_),
    .C(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__a22oi_4 _30899_ (.A1(_07934_),
    .A2(_05174_),
    .B1(_07758_),
    .B2(_05493_),
    .Y(_08559_));
 sky130_fd_sc_hd__and4_2 _30900_ (.A(_07978_),
    .B(_08174_),
    .C(_05268_),
    .D(_19920_),
    .X(_08560_));
 sky130_fd_sc_hd__nand2_2 _30901_ (.A(_19627_),
    .B(_05637_),
    .Y(_08561_));
 sky130_vsdinv _30902_ (.A(_08561_),
    .Y(_08562_));
 sky130_fd_sc_hd__o21ai_2 _30903_ (.A1(_08559_),
    .A2(_08560_),
    .B1(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__nand2_1 _30904_ (.A(_07486_),
    .B(_05236_),
    .Y(_08564_));
 sky130_fd_sc_hd__clkbuf_8 _30905_ (.A(_08174_),
    .X(_08565_));
 sky130_fd_sc_hd__nand3b_4 _30906_ (.A_N(_08564_),
    .B(_08565_),
    .C(_06073_),
    .Y(_08566_));
 sky130_fd_sc_hd__buf_8 _30907_ (.A(_07258_),
    .X(_08567_));
 sky130_fd_sc_hd__a22o_1 _30908_ (.A1(_07757_),
    .A2(_05174_),
    .B1(_08567_),
    .B2(_05378_),
    .X(_08568_));
 sky130_fd_sc_hd__nand3_2 _30909_ (.A(_08566_),
    .B(_08568_),
    .C(_08561_),
    .Y(_08569_));
 sky130_fd_sc_hd__nand2_4 _30910_ (.A(_08563_),
    .B(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__a21o_1 _30911_ (.A1(_08554_),
    .A2(_08558_),
    .B1(_08570_),
    .X(_08571_));
 sky130_fd_sc_hd__nand3_4 _30912_ (.A(_08554_),
    .B(_08558_),
    .C(_08570_),
    .Y(_08572_));
 sky130_fd_sc_hd__nand3_4 _30913_ (.A(_08537_),
    .B(_08571_),
    .C(_08572_),
    .Y(_08573_));
 sky130_fd_sc_hd__a21boi_1 _30914_ (.A1(_08169_),
    .A2(_08179_),
    .B1_N(_08165_),
    .Y(_08574_));
 sky130_fd_sc_hd__nand2_1 _30915_ (.A(_08571_),
    .B(_08572_),
    .Y(_08575_));
 sky130_fd_sc_hd__nand2_2 _30916_ (.A(_08574_),
    .B(_08575_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand2_1 _30917_ (.A(_08573_),
    .B(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__clkinv_8 _30918_ (.A(_19602_),
    .Y(_08578_));
 sky130_fd_sc_hd__buf_8 _30919_ (.A(_08578_),
    .X(_08579_));
 sky130_fd_sc_hd__buf_6 _30920_ (.A(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__nor2_2 _30921_ (.A(_08580_),
    .B(_04842_),
    .Y(_08581_));
 sky130_vsdinv _30922_ (.A(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__nand2_1 _30923_ (.A(_08577_),
    .B(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__nand3_4 _30924_ (.A(_08573_),
    .B(_08576_),
    .C(_08581_),
    .Y(_08584_));
 sky130_fd_sc_hd__nand2_2 _30925_ (.A(_08583_),
    .B(_08584_),
    .Y(_08585_));
 sky130_vsdinv _30926_ (.A(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__a22oi_4 _30927_ (.A1(_06398_),
    .A2(_06286_),
    .B1(_06838_),
    .B2(_06640_),
    .Y(_08587_));
 sky130_fd_sc_hd__nand2_1 _30928_ (.A(_06156_),
    .B(_06780_),
    .Y(_08588_));
 sky130_fd_sc_hd__nand3b_2 _30929_ (.A_N(_08588_),
    .B(_06336_),
    .C(net435),
    .Y(_08589_));
 sky130_fd_sc_hd__nand2_1 _30930_ (.A(_05731_),
    .B(_07059_),
    .Y(_08590_));
 sky130_vsdinv _30931_ (.A(_08590_),
    .Y(_08591_));
 sky130_fd_sc_hd__nand2_1 _30932_ (.A(_08589_),
    .B(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__and4_1 _30933_ (.A(_06883_),
    .B(_06019_),
    .C(_19888_),
    .D(_07281_),
    .X(_08593_));
 sky130_fd_sc_hd__o21ai_1 _30934_ (.A1(_08587_),
    .A2(_08593_),
    .B1(_08590_),
    .Y(_08594_));
 sky130_fd_sc_hd__o21a_2 _30935_ (.A1(_08587_),
    .A2(_08592_),
    .B1(_08594_),
    .X(_08595_));
 sky130_fd_sc_hd__o21ai_4 _30936_ (.A1(_08221_),
    .A2(_08218_),
    .B1(_08224_),
    .Y(_08596_));
 sky130_fd_sc_hd__buf_4 _30937_ (.A(_08219_),
    .X(_08597_));
 sky130_fd_sc_hd__a22oi_4 _30938_ (.A1(_08597_),
    .A2(_05799_),
    .B1(_06169_),
    .B2(_06119_),
    .Y(_08598_));
 sky130_fd_sc_hd__nand2_2 _30939_ (.A(_08219_),
    .B(_05798_),
    .Y(_08599_));
 sky130_fd_sc_hd__nand2_2 _30940_ (.A(_06906_),
    .B(_06118_),
    .Y(_08600_));
 sky130_fd_sc_hd__nor2_4 _30941_ (.A(_08599_),
    .B(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__nand2_2 _30942_ (.A(_06419_),
    .B(_06652_),
    .Y(_08602_));
 sky130_vsdinv _30943_ (.A(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__o21ai_2 _30944_ (.A1(_08598_),
    .A2(_08601_),
    .B1(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand2_2 _30945_ (.A(_08599_),
    .B(_08600_),
    .Y(_08605_));
 sky130_fd_sc_hd__nand3b_2 _30946_ (.A_N(_08601_),
    .B(_08602_),
    .C(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__nand3b_4 _30947_ (.A_N(_08596_),
    .B(_08604_),
    .C(_08606_),
    .Y(_08607_));
 sky130_fd_sc_hd__nand3b_4 _30948_ (.A_N(_08601_),
    .B(_08603_),
    .C(_08605_),
    .Y(_08608_));
 sky130_fd_sc_hd__o21ai_2 _30949_ (.A1(_08598_),
    .A2(_08601_),
    .B1(_08602_),
    .Y(_08609_));
 sky130_fd_sc_hd__nand3_4 _30950_ (.A(_08608_),
    .B(_08596_),
    .C(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__nand3_2 _30951_ (.A(_08595_),
    .B(_08607_),
    .C(_08610_),
    .Y(_08611_));
 sky130_vsdinv _30952_ (.A(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__a21oi_4 _30953_ (.A1(_08607_),
    .A2(_08610_),
    .B1(_08595_),
    .Y(_08613_));
 sky130_fd_sc_hd__nand2_1 _30954_ (.A(_08202_),
    .B(_08210_),
    .Y(_08614_));
 sky130_fd_sc_hd__buf_6 _30955_ (.A(_06986_),
    .X(_08615_));
 sky130_fd_sc_hd__buf_8 _30956_ (.A(_06988_),
    .X(_08616_));
 sky130_fd_sc_hd__a22oi_4 _30957_ (.A1(_08615_),
    .A2(_05770_),
    .B1(_08616_),
    .B2(_06686_),
    .Y(_08617_));
 sky130_fd_sc_hd__nand3_4 _30958_ (.A(_08190_),
    .B(_07428_),
    .C(_05481_),
    .Y(_08618_));
 sky130_fd_sc_hd__nor2_4 _30959_ (.A(net449),
    .B(_08618_),
    .Y(_08619_));
 sky130_fd_sc_hd__nand2_2 _30960_ (.A(_06992_),
    .B(_05796_),
    .Y(_08620_));
 sky130_fd_sc_hd__o21ai_2 _30961_ (.A1(_08617_),
    .A2(_08619_),
    .B1(_08620_),
    .Y(_08621_));
 sky130_vsdinv _30962_ (.A(_08620_),
    .Y(_08622_));
 sky130_fd_sc_hd__buf_6 _30963_ (.A(_08192_),
    .X(_08623_));
 sky130_fd_sc_hd__a22o_2 _30964_ (.A1(_06924_),
    .A2(_05489_),
    .B1(_08623_),
    .B2(_05958_),
    .X(_08624_));
 sky130_fd_sc_hd__o211ai_2 _30965_ (.A1(_08189_),
    .A2(_08618_),
    .B1(_08622_),
    .C1(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__o22ai_4 _30966_ (.A1(_07426_),
    .A2(_08175_),
    .B1(_08170_),
    .B2(_08173_),
    .Y(_08626_));
 sky130_fd_sc_hd__nand3_4 _30967_ (.A(_08621_),
    .B(_08625_),
    .C(_08626_),
    .Y(_08627_));
 sky130_fd_sc_hd__o21ai_2 _30968_ (.A1(_08617_),
    .A2(_08619_),
    .B1(_08622_),
    .Y(_08628_));
 sky130_fd_sc_hd__o22a_1 _30969_ (.A1(_07426_),
    .A2(_08175_),
    .B1(_08170_),
    .B2(_08173_),
    .X(_08629_));
 sky130_fd_sc_hd__o211ai_4 _30970_ (.A1(_08189_),
    .A2(_08618_),
    .B1(_08620_),
    .C1(_08624_),
    .Y(_08630_));
 sky130_fd_sc_hd__nand3_4 _30971_ (.A(_08628_),
    .B(_08629_),
    .C(_08630_),
    .Y(_08631_));
 sky130_fd_sc_hd__nor2_4 _30972_ (.A(_08200_),
    .B(_08194_),
    .Y(_08632_));
 sky130_fd_sc_hd__o2bb2ai_4 _30973_ (.A1_N(_08627_),
    .A2_N(_08631_),
    .B1(_08191_),
    .B2(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__nor2_2 _30974_ (.A(_08191_),
    .B(_08632_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand3_4 _30975_ (.A(_08631_),
    .B(_08627_),
    .C(_08634_),
    .Y(_08635_));
 sky130_fd_sc_hd__a22oi_4 _30976_ (.A1(_08207_),
    .A2(_08614_),
    .B1(_08633_),
    .B2(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__and3_1 _30977_ (.A(_08195_),
    .B(_08196_),
    .C(_08201_),
    .X(_08637_));
 sky130_fd_sc_hd__a31oi_2 _30978_ (.A1(_08203_),
    .A2(_08205_),
    .A3(_08206_),
    .B1(_08210_),
    .Y(_08638_));
 sky130_fd_sc_hd__o211a_4 _30979_ (.A1(_08637_),
    .A2(_08638_),
    .B1(_08635_),
    .C1(_08633_),
    .X(_08639_));
 sky130_fd_sc_hd__o22ai_4 _30980_ (.A1(_08612_),
    .A2(_08613_),
    .B1(_08636_),
    .B2(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__nand2_1 _30981_ (.A(_08207_),
    .B(_08211_),
    .Y(_08641_));
 sky130_fd_sc_hd__nand2_2 _30982_ (.A(_08641_),
    .B(_08202_),
    .Y(_08642_));
 sky130_fd_sc_hd__a21o_1 _30983_ (.A1(_08633_),
    .A2(_08635_),
    .B1(_08642_),
    .X(_08643_));
 sky130_fd_sc_hd__o211a_1 _30984_ (.A1(_08587_),
    .A2(_08592_),
    .B1(_08594_),
    .C1(_08610_),
    .X(_08644_));
 sky130_fd_sc_hd__a21oi_4 _30985_ (.A1(_08644_),
    .A2(_08607_),
    .B1(_08613_),
    .Y(_08645_));
 sky130_fd_sc_hd__nand3_4 _30986_ (.A(_08642_),
    .B(_08633_),
    .C(_08635_),
    .Y(_08646_));
 sky130_fd_sc_hd__nand3_2 _30987_ (.A(_08643_),
    .B(_08645_),
    .C(_08646_),
    .Y(_08647_));
 sky130_fd_sc_hd__nand3_4 _30988_ (.A(_08640_),
    .B(_08184_),
    .C(_08647_),
    .Y(_08648_));
 sky130_fd_sc_hd__o21ai_2 _30989_ (.A1(_08636_),
    .A2(_08639_),
    .B1(_08645_),
    .Y(_08649_));
 sky130_fd_sc_hd__nand3_2 _30990_ (.A(_08185_),
    .B(_08181_),
    .C(_08182_),
    .Y(_08650_));
 sky130_fd_sc_hd__a21o_1 _30991_ (.A1(_08607_),
    .A2(_08610_),
    .B1(_08595_),
    .X(_08651_));
 sky130_fd_sc_hd__nand2_2 _30992_ (.A(_08651_),
    .B(_08611_),
    .Y(_08652_));
 sky130_fd_sc_hd__nand3_2 _30993_ (.A(_08643_),
    .B(_08646_),
    .C(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__nand3_4 _30994_ (.A(_08649_),
    .B(_08650_),
    .C(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__nor2_8 _30995_ (.A(_08252_),
    .B(_08216_),
    .Y(_08655_));
 sky130_fd_sc_hd__o2bb2ai_2 _30996_ (.A1_N(_08648_),
    .A2_N(_08654_),
    .B1(_08214_),
    .B2(_08655_),
    .Y(_08656_));
 sky130_fd_sc_hd__nor2_8 _30997_ (.A(_08214_),
    .B(_08655_),
    .Y(_08657_));
 sky130_fd_sc_hd__nand3_4 _30998_ (.A(_08654_),
    .B(_08648_),
    .C(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand3_4 _30999_ (.A(_08586_),
    .B(_08656_),
    .C(_08658_),
    .Y(_08659_));
 sky130_fd_sc_hd__nand2_1 _31000_ (.A(_08656_),
    .B(_08658_),
    .Y(_08660_));
 sky130_fd_sc_hd__a21oi_1 _31001_ (.A1(_08660_),
    .A2(_08585_),
    .B1(_08272_),
    .Y(_08661_));
 sky130_vsdinv _31002_ (.A(_08583_),
    .Y(_08662_));
 sky130_vsdinv _31003_ (.A(_08584_),
    .Y(_08663_));
 sky130_fd_sc_hd__a2bb2oi_4 _31004_ (.A1_N(_08214_),
    .A2_N(_08655_),
    .B1(_08648_),
    .B2(_08654_),
    .Y(_08664_));
 sky130_fd_sc_hd__nor2_1 _31005_ (.A(_08214_),
    .B(_08246_),
    .Y(_08665_));
 sky130_fd_sc_hd__o211a_2 _31006_ (.A1(_08216_),
    .A2(_08665_),
    .B1(_08648_),
    .C1(_08654_),
    .X(_08666_));
 sky130_fd_sc_hd__o22ai_4 _31007_ (.A1(_08662_),
    .A2(_08663_),
    .B1(_08664_),
    .B2(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__a22oi_2 _31008_ (.A1(_08390_),
    .A2(_08271_),
    .B1(_08667_),
    .B2(_08659_),
    .Y(_08668_));
 sky130_fd_sc_hd__a21oi_2 _31009_ (.A1(_08659_),
    .A2(_08661_),
    .B1(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__o21ai_4 _31010_ (.A1(_08533_),
    .A2(_08535_),
    .B1(_08669_),
    .Y(_08670_));
 sky130_fd_sc_hd__a21oi_2 _31011_ (.A1(_08656_),
    .A2(_08658_),
    .B1(_08586_),
    .Y(_08671_));
 sky130_fd_sc_hd__nor3_4 _31012_ (.A(_08585_),
    .B(_08664_),
    .C(_08666_),
    .Y(_08672_));
 sky130_fd_sc_hd__o22ai_4 _31013_ (.A1(_08265_),
    .A2(_08277_),
    .B1(_08671_),
    .B2(_08672_),
    .Y(_08673_));
 sky130_fd_sc_hd__nand3_4 _31014_ (.A(_08383_),
    .B(_08667_),
    .C(_08659_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand2_2 _31015_ (.A(_08673_),
    .B(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__nand2_4 _31016_ (.A(_08534_),
    .B(_08531_),
    .Y(_08676_));
 sky130_fd_sc_hd__nand3_4 _31017_ (.A(_08532_),
    .B(_08524_),
    .C(_08530_),
    .Y(_08677_));
 sky130_fd_sc_hd__nand3_4 _31018_ (.A(_08675_),
    .B(_08676_),
    .C(_08677_),
    .Y(_08678_));
 sky130_fd_sc_hd__nand3_4 _31019_ (.A(_08440_),
    .B(_08670_),
    .C(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__nand3_1 _31020_ (.A(_08387_),
    .B(_08386_),
    .C(_08385_),
    .Y(_08680_));
 sky130_fd_sc_hd__nand2_1 _31021_ (.A(_08680_),
    .B(_08391_),
    .Y(_08681_));
 sky130_fd_sc_hd__o21ai_2 _31022_ (.A1(_08533_),
    .A2(_08535_),
    .B1(_08675_),
    .Y(_08682_));
 sky130_vsdinv _31023_ (.A(_08530_),
    .Y(_08683_));
 sky130_fd_sc_hd__nand2_2 _31024_ (.A(_08532_),
    .B(_08524_),
    .Y(_08684_));
 sky130_fd_sc_hd__o2111ai_4 _31025_ (.A1(_08683_),
    .A2(_08684_),
    .B1(_08674_),
    .C1(_08673_),
    .D1(_08676_),
    .Y(_08685_));
 sky130_fd_sc_hd__nand3_4 _31026_ (.A(_08681_),
    .B(_08682_),
    .C(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand2_1 _31027_ (.A(_08679_),
    .B(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__nand2_1 _31028_ (.A(_08385_),
    .B(_08374_),
    .Y(_08688_));
 sky130_fd_sc_hd__nand2_1 _31029_ (.A(_08361_),
    .B(_08357_),
    .Y(_08689_));
 sky130_fd_sc_hd__nand2_2 _31030_ (.A(_08688_),
    .B(_08689_),
    .Y(_08690_));
 sky130_vsdinv _31031_ (.A(_08689_),
    .Y(_08691_));
 sky130_fd_sc_hd__nand3_2 _31032_ (.A(_08385_),
    .B(_08374_),
    .C(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__nand2_2 _31033_ (.A(_08690_),
    .B(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__nand2_1 _31034_ (.A(_08687_),
    .B(_08693_),
    .Y(_08694_));
 sky130_fd_sc_hd__nand2_1 _31035_ (.A(_08395_),
    .B(_08414_),
    .Y(_08695_));
 sky130_fd_sc_hd__nand2_1 _31036_ (.A(_08695_),
    .B(_08389_),
    .Y(_08696_));
 sky130_fd_sc_hd__and2_2 _31037_ (.A(_08690_),
    .B(_08692_),
    .X(_08697_));
 sky130_fd_sc_hd__nand3_4 _31038_ (.A(_08679_),
    .B(_08686_),
    .C(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__nand3_4 _31039_ (.A(_08694_),
    .B(_08696_),
    .C(_08698_),
    .Y(_08699_));
 sky130_vsdinv _31040_ (.A(_08688_),
    .Y(_08700_));
 sky130_fd_sc_hd__nor2_1 _31041_ (.A(_08689_),
    .B(_08700_),
    .Y(_08701_));
 sky130_fd_sc_hd__nor2_1 _31042_ (.A(_08691_),
    .B(_08688_),
    .Y(_08702_));
 sky130_fd_sc_hd__o2bb2ai_2 _31043_ (.A1_N(_08686_),
    .A2_N(_08679_),
    .B1(_08701_),
    .B2(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__a21boi_4 _31044_ (.A1(_08395_),
    .A2(_08414_),
    .B1_N(_08389_),
    .Y(_08704_));
 sky130_fd_sc_hd__nand3_2 _31045_ (.A(_08679_),
    .B(_08686_),
    .C(_08693_),
    .Y(_08705_));
 sky130_fd_sc_hd__nand3_4 _31046_ (.A(_08703_),
    .B(_08704_),
    .C(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__nand2_1 _31047_ (.A(_08699_),
    .B(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__nand2_1 _31048_ (.A(_08707_),
    .B(_08411_),
    .Y(_08708_));
 sky130_fd_sc_hd__a21boi_4 _31049_ (.A1(_08410_),
    .A2(_07890_),
    .B1_N(_08417_),
    .Y(_08709_));
 sky130_fd_sc_hd__nand3_2 _31050_ (.A(_08699_),
    .B(_08706_),
    .C(_08406_),
    .Y(_08710_));
 sky130_fd_sc_hd__nand3_4 _31051_ (.A(_08708_),
    .B(_08709_),
    .C(_08710_),
    .Y(_08711_));
 sky130_fd_sc_hd__nand2_1 _31052_ (.A(_08707_),
    .B(_08406_),
    .Y(_08712_));
 sky130_fd_sc_hd__nand2_1 _31053_ (.A(_08410_),
    .B(_07890_),
    .Y(_08713_));
 sky130_fd_sc_hd__nand2_2 _31054_ (.A(_08713_),
    .B(_08417_),
    .Y(_08714_));
 sky130_fd_sc_hd__nand3_2 _31055_ (.A(_08699_),
    .B(_08706_),
    .C(_08411_),
    .Y(_08715_));
 sky130_fd_sc_hd__nand3_4 _31056_ (.A(_08712_),
    .B(_08714_),
    .C(_08715_),
    .Y(_08716_));
 sky130_fd_sc_hd__nand2_4 _31057_ (.A(_08711_),
    .B(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__nor2_2 _31058_ (.A(_08428_),
    .B(_08142_),
    .Y(_08718_));
 sky130_fd_sc_hd__nand3_2 _31059_ (.A(_08718_),
    .B(_07633_),
    .C(_07884_),
    .Y(_08719_));
 sky130_vsdinv _31060_ (.A(_08422_),
    .Y(_08720_));
 sky130_fd_sc_hd__o21ai_1 _31061_ (.A1(_08141_),
    .A2(_08720_),
    .B1(_08427_),
    .Y(_08721_));
 sky130_fd_sc_hd__a21oi_2 _31062_ (.A1(_08718_),
    .A2(_08144_),
    .B1(_08721_),
    .Y(_08722_));
 sky130_fd_sc_hd__o21ai_4 _31063_ (.A1(_08719_),
    .A2(_07638_),
    .B1(_08722_),
    .Y(_08723_));
 sky130_vsdinv _31064_ (.A(_08723_),
    .Y(_08724_));
 sky130_fd_sc_hd__and3_1 _31065_ (.A(_08439_),
    .B(_08717_),
    .C(_08724_),
    .X(_08725_));
 sky130_fd_sc_hd__and2_1 _31066_ (.A(_08439_),
    .B(_08724_),
    .X(_08726_));
 sky130_fd_sc_hd__nor2_2 _31067_ (.A(_08717_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__nor2_4 _31068_ (.A(_08725_),
    .B(_08727_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand3_1 _31069_ (.A(_08676_),
    .B(_08673_),
    .C(_08677_),
    .Y(_08728_));
 sky130_fd_sc_hd__nand2_2 _31070_ (.A(_08728_),
    .B(_08674_),
    .Y(_08729_));
 sky130_vsdinv _31071_ (.A(_08464_),
    .Y(_08730_));
 sky130_fd_sc_hd__nand3_4 _31072_ (.A(_05591_),
    .B(_05842_),
    .C(_07345_),
    .Y(_08731_));
 sky130_fd_sc_hd__nor2_4 _31073_ (.A(net470),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__nand2_2 _31074_ (.A(_05259_),
    .B(_07556_),
    .Y(_08733_));
 sky130_fd_sc_hd__buf_6 _31075_ (.A(_07050_),
    .X(_08734_));
 sky130_fd_sc_hd__buf_6 _31076_ (.A(_07554_),
    .X(_08735_));
 sky130_fd_sc_hd__a22o_2 _31077_ (.A1(_05837_),
    .A2(_08734_),
    .B1(_06077_),
    .B2(_08735_),
    .X(_08736_));
 sky130_fd_sc_hd__nand3b_2 _31078_ (.A_N(_08732_),
    .B(_08733_),
    .C(_08736_),
    .Y(_08737_));
 sky130_fd_sc_hd__a22o_1 _31079_ (.A1(_06156_),
    .A2(_06780_),
    .B1(_05883_),
    .B2(_07327_),
    .X(_08738_));
 sky130_fd_sc_hd__a21oi_4 _31080_ (.A1(_08738_),
    .A2(_08591_),
    .B1(_08593_),
    .Y(_08739_));
 sky130_fd_sc_hd__a22oi_4 _31081_ (.A1(_06502_),
    .A2(_07056_),
    .B1(_06835_),
    .B2(_08735_),
    .Y(_08740_));
 sky130_vsdinv _31082_ (.A(_08733_),
    .Y(_08741_));
 sky130_fd_sc_hd__o21ai_2 _31083_ (.A1(_08740_),
    .A2(_08732_),
    .B1(_08741_),
    .Y(_08742_));
 sky130_fd_sc_hd__nand3_4 _31084_ (.A(_08737_),
    .B(_08739_),
    .C(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__o21ai_2 _31085_ (.A1(_08740_),
    .A2(_08732_),
    .B1(_08733_),
    .Y(_08744_));
 sky130_fd_sc_hd__clkbuf_2 _31086_ (.A(net470),
    .X(_08745_));
 sky130_fd_sc_hd__o211ai_2 _31087_ (.A1(net438),
    .A2(_08731_),
    .B1(_08741_),
    .C1(_08736_),
    .Y(_08746_));
 sky130_fd_sc_hd__o21ai_2 _31088_ (.A1(_08590_),
    .A2(_08587_),
    .B1(_08589_),
    .Y(_08747_));
 sky130_fd_sc_hd__nand3_4 _31089_ (.A(_08744_),
    .B(_08746_),
    .C(_08747_),
    .Y(_08748_));
 sky130_fd_sc_hd__a21oi_2 _31090_ (.A1(_08449_),
    .A2(_08448_),
    .B1(_08443_),
    .Y(_08749_));
 sky130_vsdinv _31091_ (.A(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__a21o_2 _31092_ (.A1(_08743_),
    .A2(_08748_),
    .B1(_08750_),
    .X(_08751_));
 sky130_fd_sc_hd__nand3_4 _31093_ (.A(_08743_),
    .B(_08748_),
    .C(_08750_),
    .Y(_08752_));
 sky130_vsdinv _31094_ (.A(_08609_),
    .Y(_08753_));
 sky130_fd_sc_hd__nand2_1 _31095_ (.A(_08608_),
    .B(_08596_),
    .Y(_08754_));
 sky130_fd_sc_hd__o2bb2ai_4 _31096_ (.A1_N(_08607_),
    .A2_N(_08595_),
    .B1(_08753_),
    .B2(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__a21oi_4 _31097_ (.A1(_08751_),
    .A2(_08752_),
    .B1(_08755_),
    .Y(_08756_));
 sky130_vsdinv _31098_ (.A(_08748_),
    .Y(_08757_));
 sky130_fd_sc_hd__nand2_1 _31099_ (.A(_08743_),
    .B(_08750_),
    .Y(_08758_));
 sky130_fd_sc_hd__o211a_1 _31100_ (.A1(_08757_),
    .A2(_08758_),
    .B1(_08751_),
    .C1(_08755_),
    .X(_08759_));
 sky130_fd_sc_hd__o22ai_4 _31101_ (.A1(_08465_),
    .A2(_08730_),
    .B1(_08756_),
    .B2(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__o21a_1 _31102_ (.A1(_08467_),
    .A2(_08463_),
    .B1(_08470_),
    .X(_08761_));
 sky130_fd_sc_hd__a21o_1 _31103_ (.A1(_08751_),
    .A2(_08752_),
    .B1(_08755_),
    .X(_08762_));
 sky130_fd_sc_hd__nand3_4 _31104_ (.A(_08755_),
    .B(_08751_),
    .C(_08752_),
    .Y(_08763_));
 sky130_fd_sc_hd__nor2_8 _31105_ (.A(_08465_),
    .B(_08730_),
    .Y(_08764_));
 sky130_fd_sc_hd__nand3_2 _31106_ (.A(_08762_),
    .B(_08763_),
    .C(_08764_),
    .Y(_08765_));
 sky130_fd_sc_hd__nand3_4 _31107_ (.A(_08760_),
    .B(_08761_),
    .C(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__o21ai_2 _31108_ (.A1(_08756_),
    .A2(_08759_),
    .B1(_08764_),
    .Y(_08767_));
 sky130_fd_sc_hd__o21ai_2 _31109_ (.A1(_08467_),
    .A2(_08463_),
    .B1(_08470_),
    .Y(_08768_));
 sky130_fd_sc_hd__nand3b_2 _31110_ (.A_N(_08764_),
    .B(_08762_),
    .C(_08763_),
    .Y(_08769_));
 sky130_fd_sc_hd__nand3_4 _31111_ (.A(_08767_),
    .B(_08768_),
    .C(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__nand2_2 _31112_ (.A(_08500_),
    .B(_08501_),
    .Y(_08771_));
 sky130_fd_sc_hd__nand2_1 _31113_ (.A(_08771_),
    .B(_08502_),
    .Y(_08772_));
 sky130_fd_sc_hd__clkbuf_4 _31114_ (.A(\pcpi_mul.rs1[24] ),
    .X(_08773_));
 sky130_fd_sc_hd__and4_2 _31115_ (.A(_05117_),
    .B(_05119_),
    .C(_08773_),
    .D(_19858_),
    .X(_08774_));
 sky130_fd_sc_hd__a22o_1 _31116_ (.A1(_06636_),
    .A2(_19858_),
    .B1(_05119_),
    .B2(_08773_),
    .X(_08775_));
 sky130_vsdinv _31117_ (.A(_08775_),
    .Y(_08776_));
 sky130_fd_sc_hd__nor2_2 _31118_ (.A(_05132_),
    .B(_08043_),
    .Y(_08777_));
 sky130_fd_sc_hd__o21ai_1 _31119_ (.A1(_08774_),
    .A2(_08776_),
    .B1(_08777_),
    .Y(_08778_));
 sky130_vsdinv _31120_ (.A(_08777_),
    .Y(_08779_));
 sky130_fd_sc_hd__nand3b_1 _31121_ (.A_N(_08774_),
    .B(_08779_),
    .C(_08775_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand2_1 _31122_ (.A(_08778_),
    .B(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__nand2_2 _31123_ (.A(_05211_),
    .B(_07542_),
    .Y(_08782_));
 sky130_fd_sc_hd__nand2_2 _31124_ (.A(_19672_),
    .B(_07686_),
    .Y(_08783_));
 sky130_fd_sc_hd__nor2_4 _31125_ (.A(_08782_),
    .B(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__nand2_2 _31126_ (.A(_08782_),
    .B(_08783_),
    .Y(_08785_));
 sky130_vsdinv _31127_ (.A(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__buf_4 _31128_ (.A(\pcpi_mul.rs1[25] ),
    .X(_08787_));
 sky130_fd_sc_hd__nand2_2 _31129_ (.A(_05171_),
    .B(_08787_),
    .Y(_08788_));
 sky130_vsdinv _31130_ (.A(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__o21ai_2 _31131_ (.A1(_08784_),
    .A2(_08786_),
    .B1(_08789_),
    .Y(_08790_));
 sky130_vsdinv _31132_ (.A(_08784_),
    .Y(_08791_));
 sky130_fd_sc_hd__nand3_2 _31133_ (.A(_08791_),
    .B(_08788_),
    .C(_08785_),
    .Y(_08792_));
 sky130_fd_sc_hd__a21oi_2 _31134_ (.A1(_08488_),
    .A2(_08486_),
    .B1(_08484_),
    .Y(_08793_));
 sky130_fd_sc_hd__nand3_4 _31135_ (.A(_08790_),
    .B(_08792_),
    .C(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__o21ai_2 _31136_ (.A1(_08784_),
    .A2(_08786_),
    .B1(_08788_),
    .Y(_08795_));
 sky130_fd_sc_hd__nand3_2 _31137_ (.A(_08791_),
    .B(_08789_),
    .C(_08785_),
    .Y(_08796_));
 sky130_fd_sc_hd__a21o_1 _31138_ (.A1(_08488_),
    .A2(_08486_),
    .B1(_08484_),
    .X(_08797_));
 sky130_fd_sc_hd__nand3_4 _31139_ (.A(_08795_),
    .B(_08796_),
    .C(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__nand3_2 _31140_ (.A(_08781_),
    .B(_08794_),
    .C(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__nand2_1 _31141_ (.A(_08798_),
    .B(_08794_),
    .Y(_08800_));
 sky130_fd_sc_hd__o21ai_1 _31142_ (.A1(_08774_),
    .A2(_08776_),
    .B1(_08779_),
    .Y(_08801_));
 sky130_fd_sc_hd__nand3b_2 _31143_ (.A_N(_08774_),
    .B(_08777_),
    .C(_08775_),
    .Y(_08802_));
 sky130_fd_sc_hd__nand2_1 _31144_ (.A(_08801_),
    .B(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__nand2_1 _31145_ (.A(_08800_),
    .B(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__nand3_4 _31146_ (.A(_08772_),
    .B(_08799_),
    .C(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__nand3_2 _31147_ (.A(_08803_),
    .B(_08794_),
    .C(_08798_),
    .Y(_08806_));
 sky130_fd_sc_hd__nand2_1 _31148_ (.A(_08800_),
    .B(_08781_),
    .Y(_08807_));
 sky130_fd_sc_hd__o2111ai_4 _31149_ (.A1(_08495_),
    .A2(_08494_),
    .B1(_08771_),
    .C1(_08806_),
    .D1(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__nor2_2 _31150_ (.A(_08475_),
    .B(_08478_),
    .Y(_08809_));
 sky130_fd_sc_hd__nor2_4 _31151_ (.A(_08809_),
    .B(_08483_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand3_2 _31152_ (.A(_08805_),
    .B(_08808_),
    .C(_08810_),
    .Y(_08811_));
 sky130_vsdinv _31153_ (.A(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__nand2_2 _31154_ (.A(_08805_),
    .B(_08808_),
    .Y(_08813_));
 sky130_vsdinv _31155_ (.A(_08810_),
    .Y(_08814_));
 sky130_fd_sc_hd__and2_1 _31156_ (.A(_08813_),
    .B(_08814_),
    .X(_08815_));
 sky130_fd_sc_hd__o2bb2ai_2 _31157_ (.A1_N(_08766_),
    .A2_N(_08770_),
    .B1(_08812_),
    .B2(_08815_),
    .Y(_08816_));
 sky130_fd_sc_hd__a21boi_4 _31158_ (.A1(_08654_),
    .A2(_08657_),
    .B1_N(_08648_),
    .Y(_08817_));
 sky130_fd_sc_hd__nand2_1 _31159_ (.A(_08808_),
    .B(_08814_),
    .Y(_08818_));
 sky130_vsdinv _31160_ (.A(_08805_),
    .Y(_08819_));
 sky130_fd_sc_hd__nand2_1 _31161_ (.A(_08813_),
    .B(_08810_),
    .Y(_08820_));
 sky130_fd_sc_hd__o21ai_1 _31162_ (.A1(_08818_),
    .A2(_08819_),
    .B1(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__nand3_2 _31163_ (.A(_08821_),
    .B(_08770_),
    .C(_08766_),
    .Y(_08822_));
 sky130_fd_sc_hd__nand3_4 _31164_ (.A(_08816_),
    .B(_08817_),
    .C(_08822_),
    .Y(_08823_));
 sky130_fd_sc_hd__nor2_1 _31165_ (.A(_08810_),
    .B(_08813_),
    .Y(_08824_));
 sky130_fd_sc_hd__and2_1 _31166_ (.A(_08813_),
    .B(_08810_),
    .X(_08825_));
 sky130_fd_sc_hd__o2bb2ai_2 _31167_ (.A1_N(_08766_),
    .A2_N(_08770_),
    .B1(_08824_),
    .B2(_08825_),
    .Y(_08826_));
 sky130_fd_sc_hd__nand2_1 _31168_ (.A(_08654_),
    .B(_08657_),
    .Y(_08827_));
 sky130_fd_sc_hd__nand2_2 _31169_ (.A(_08827_),
    .B(_08648_),
    .Y(_08828_));
 sky130_fd_sc_hd__nand2_1 _31170_ (.A(_08813_),
    .B(_08814_),
    .Y(_08829_));
 sky130_fd_sc_hd__nand2_2 _31171_ (.A(_08829_),
    .B(_08811_),
    .Y(_08830_));
 sky130_fd_sc_hd__nand3_4 _31172_ (.A(_08830_),
    .B(_08770_),
    .C(_08766_),
    .Y(_08831_));
 sky130_fd_sc_hd__nand3_4 _31173_ (.A(_08826_),
    .B(_08828_),
    .C(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__nor2_2 _31174_ (.A(_08474_),
    .B(_08512_),
    .Y(_08833_));
 sky130_fd_sc_hd__o2bb2ai_4 _31175_ (.A1_N(_08823_),
    .A2_N(_08832_),
    .B1(_08472_),
    .B2(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__o21ai_4 _31176_ (.A1(_08472_),
    .A2(_08522_),
    .B1(_08518_),
    .Y(_08835_));
 sky130_fd_sc_hd__nand3_4 _31177_ (.A(_08823_),
    .B(_08832_),
    .C(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__nand2_1 _31178_ (.A(_08834_),
    .B(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__nor2_4 _31179_ (.A(_08645_),
    .B(_08639_),
    .Y(_08838_));
 sky130_fd_sc_hd__o21ai_1 _31180_ (.A1(_08599_),
    .A2(_08600_),
    .B1(_08602_),
    .Y(_08839_));
 sky130_fd_sc_hd__nand2_2 _31181_ (.A(_08839_),
    .B(_08605_),
    .Y(_08840_));
 sky130_fd_sc_hd__a22oi_4 _31182_ (.A1(_06341_),
    .A2(_19898_),
    .B1(_06416_),
    .B2(_19894_),
    .Y(_08841_));
 sky130_fd_sc_hd__and4_2 _31183_ (.A(_08219_),
    .B(_06906_),
    .C(_07502_),
    .D(_06657_),
    .X(_08842_));
 sky130_fd_sc_hd__nand2_2 _31184_ (.A(_19649_),
    .B(_06779_),
    .Y(_08843_));
 sky130_fd_sc_hd__o21ai_2 _31185_ (.A1(_08841_),
    .A2(_08842_),
    .B1(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__nand2_1 _31186_ (.A(_07007_),
    .B(_06118_),
    .Y(_08845_));
 sky130_fd_sc_hd__nand3b_4 _31187_ (.A_N(_08845_),
    .B(_06422_),
    .C(_06650_),
    .Y(_08846_));
 sky130_vsdinv _31188_ (.A(_08843_),
    .Y(_08847_));
 sky130_fd_sc_hd__a22o_2 _31189_ (.A1(_06414_),
    .A2(_06440_),
    .B1(_06345_),
    .B2(_06652_),
    .X(_08848_));
 sky130_fd_sc_hd__nand3_2 _31190_ (.A(_08846_),
    .B(_08847_),
    .C(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__nand3b_4 _31191_ (.A_N(_08840_),
    .B(_08844_),
    .C(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__o21ai_2 _31192_ (.A1(_08841_),
    .A2(_08842_),
    .B1(_08847_),
    .Y(_08851_));
 sky130_fd_sc_hd__nand3_2 _31193_ (.A(_08846_),
    .B(_08843_),
    .C(_08848_),
    .Y(_08852_));
 sky130_fd_sc_hd__nand3_4 _31194_ (.A(_08851_),
    .B(_08852_),
    .C(_08840_),
    .Y(_08853_));
 sky130_fd_sc_hd__a22oi_4 _31195_ (.A1(_06018_),
    .A2(_07330_),
    .B1(_06335_),
    .B2(_19884_),
    .Y(_08854_));
 sky130_fd_sc_hd__nand2_2 _31196_ (.A(_06017_),
    .B(_06808_),
    .Y(_08855_));
 sky130_fd_sc_hd__nand2_1 _31197_ (.A(_05882_),
    .B(_07322_),
    .Y(_08856_));
 sky130_fd_sc_hd__nor2_1 _31198_ (.A(_08855_),
    .B(_08856_),
    .Y(_08857_));
 sky130_fd_sc_hd__nand2_2 _31199_ (.A(_06013_),
    .B(_06654_),
    .Y(_08858_));
 sky130_fd_sc_hd__o21bai_2 _31200_ (.A1(_08854_),
    .A2(_08857_),
    .B1_N(_08858_),
    .Y(_08859_));
 sky130_fd_sc_hd__nand3b_4 _31201_ (.A_N(_08855_),
    .B(_06159_),
    .C(_07323_),
    .Y(_08860_));
 sky130_fd_sc_hd__nand2_1 _31202_ (.A(_08855_),
    .B(_08856_),
    .Y(_08861_));
 sky130_fd_sc_hd__nand3_2 _31203_ (.A(_08860_),
    .B(_08858_),
    .C(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__nand2_4 _31204_ (.A(_08859_),
    .B(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__nand3_2 _31205_ (.A(_08850_),
    .B(_08853_),
    .C(_08863_),
    .Y(_08864_));
 sky130_vsdinv _31206_ (.A(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__a21oi_4 _31207_ (.A1(_08850_),
    .A2(_08853_),
    .B1(_08863_),
    .Y(_08866_));
 sky130_fd_sc_hd__nand3_4 _31208_ (.A(_07923_),
    .B(_08192_),
    .C(_19906_),
    .Y(_08867_));
 sky130_fd_sc_hd__nor2_8 _31209_ (.A(_05802_),
    .B(_08867_),
    .Y(_08868_));
 sky130_fd_sc_hd__nand2_2 _31210_ (.A(_06992_),
    .B(_05643_),
    .Y(_08869_));
 sky130_fd_sc_hd__a22o_2 _31211_ (.A1(_07744_),
    .A2(_05661_),
    .B1(_07928_),
    .B2(_06494_),
    .X(_08870_));
 sky130_fd_sc_hd__nand3b_2 _31212_ (.A_N(_08868_),
    .B(_08869_),
    .C(_08870_),
    .Y(_08871_));
 sky130_fd_sc_hd__a21oi_4 _31213_ (.A1(_08568_),
    .A2(_08562_),
    .B1(_08560_),
    .Y(_08872_));
 sky130_fd_sc_hd__buf_6 _31214_ (.A(_06988_),
    .X(_08873_));
 sky130_fd_sc_hd__a22oi_4 _31215_ (.A1(_06924_),
    .A2(_19907_),
    .B1(_08873_),
    .B2(_06257_),
    .Y(_08874_));
 sky130_vsdinv _31216_ (.A(_08869_),
    .Y(_08875_));
 sky130_fd_sc_hd__o21ai_2 _31217_ (.A1(_08874_),
    .A2(_08868_),
    .B1(_08875_),
    .Y(_08876_));
 sky130_fd_sc_hd__nand3_4 _31218_ (.A(_08871_),
    .B(_08872_),
    .C(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__o21ai_2 _31219_ (.A1(_08874_),
    .A2(_08868_),
    .B1(_08869_),
    .Y(_08878_));
 sky130_fd_sc_hd__o21ai_2 _31220_ (.A1(_08561_),
    .A2(_08559_),
    .B1(_08566_),
    .Y(_08879_));
 sky130_fd_sc_hd__o211ai_2 _31221_ (.A1(_05803_),
    .A2(_08867_),
    .B1(_08875_),
    .C1(_08870_),
    .Y(_08880_));
 sky130_fd_sc_hd__nand3_4 _31222_ (.A(_08878_),
    .B(_08879_),
    .C(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__a21oi_4 _31223_ (.A1(_08624_),
    .A2(_08622_),
    .B1(_08619_),
    .Y(_08882_));
 sky130_vsdinv _31224_ (.A(_08882_),
    .Y(_08883_));
 sky130_fd_sc_hd__a21o_2 _31225_ (.A1(_08877_),
    .A2(_08881_),
    .B1(_08883_),
    .X(_08884_));
 sky130_fd_sc_hd__nand3_4 _31226_ (.A(_08877_),
    .B(_08881_),
    .C(_08883_),
    .Y(_08885_));
 sky130_fd_sc_hd__nand2_1 _31227_ (.A(_08631_),
    .B(_08634_),
    .Y(_08886_));
 sky130_fd_sc_hd__nand2_4 _31228_ (.A(_08886_),
    .B(_08627_),
    .Y(_08887_));
 sky130_fd_sc_hd__a21oi_4 _31229_ (.A1(_08884_),
    .A2(_08885_),
    .B1(_08887_),
    .Y(_08888_));
 sky130_vsdinv _31230_ (.A(_08881_),
    .Y(_08889_));
 sky130_fd_sc_hd__nand2_1 _31231_ (.A(_08877_),
    .B(_08883_),
    .Y(_08890_));
 sky130_fd_sc_hd__o211a_2 _31232_ (.A1(_08889_),
    .A2(_08890_),
    .B1(_08887_),
    .C1(_08884_),
    .X(_08891_));
 sky130_fd_sc_hd__o22ai_4 _31233_ (.A1(_08865_),
    .A2(_08866_),
    .B1(_08888_),
    .B2(_08891_),
    .Y(_08892_));
 sky130_vsdinv _31234_ (.A(_08573_),
    .Y(_08893_));
 sky130_fd_sc_hd__a21o_1 _31235_ (.A1(_08884_),
    .A2(_08885_),
    .B1(_08887_),
    .X(_08894_));
 sky130_fd_sc_hd__nand3_4 _31236_ (.A(_08884_),
    .B(_08887_),
    .C(_08885_),
    .Y(_08895_));
 sky130_fd_sc_hd__nor2_4 _31237_ (.A(_08866_),
    .B(_08865_),
    .Y(_08896_));
 sky130_fd_sc_hd__nand3_2 _31238_ (.A(_08894_),
    .B(_08895_),
    .C(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__nand3_4 _31239_ (.A(_08892_),
    .B(_08893_),
    .C(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__o21ai_4 _31240_ (.A1(_08888_),
    .A2(_08891_),
    .B1(_08896_),
    .Y(_08899_));
 sky130_fd_sc_hd__a21o_1 _31241_ (.A1(_08850_),
    .A2(_08853_),
    .B1(_08863_),
    .X(_08900_));
 sky130_fd_sc_hd__nand2_2 _31242_ (.A(_08900_),
    .B(_08864_),
    .Y(_08901_));
 sky130_fd_sc_hd__nand3_4 _31243_ (.A(_08894_),
    .B(_08895_),
    .C(_08901_),
    .Y(_08902_));
 sky130_fd_sc_hd__nand3_4 _31244_ (.A(_08899_),
    .B(_08573_),
    .C(_08902_),
    .Y(_08903_));
 sky130_fd_sc_hd__a2bb2oi_4 _31245_ (.A1_N(_08636_),
    .A2_N(_08838_),
    .B1(_08898_),
    .B2(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__nor2_2 _31246_ (.A(_08652_),
    .B(_08636_),
    .Y(_08905_));
 sky130_fd_sc_hd__o211a_1 _31247_ (.A1(_08639_),
    .A2(_08905_),
    .B1(_08898_),
    .C1(_08903_),
    .X(_08906_));
 sky130_fd_sc_hd__nand2_2 _31248_ (.A(_08572_),
    .B(_08554_),
    .Y(_08907_));
 sky130_fd_sc_hd__buf_8 _31249_ (.A(_08539_),
    .X(_08908_));
 sky130_fd_sc_hd__a22oi_4 _31250_ (.A1(_08908_),
    .A2(_06020_),
    .B1(_08550_),
    .B2(_05264_),
    .Y(_08909_));
 sky130_fd_sc_hd__nand2_2 _31251_ (.A(_08539_),
    .B(_07828_),
    .Y(_08910_));
 sky130_fd_sc_hd__nand2_2 _31252_ (.A(_08154_),
    .B(_05695_),
    .Y(_08911_));
 sky130_fd_sc_hd__nor2_4 _31253_ (.A(_08910_),
    .B(_08911_),
    .Y(_08912_));
 sky130_fd_sc_hd__nand2_2 _31254_ (.A(_19615_),
    .B(_05173_),
    .Y(_08913_));
 sky130_vsdinv _31255_ (.A(_08913_),
    .Y(_08914_));
 sky130_fd_sc_hd__o21ai_2 _31256_ (.A1(_08909_),
    .A2(_08912_),
    .B1(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__nand3b_4 _31257_ (.A_N(_08910_),
    .B(_08541_),
    .C(_05838_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand2_2 _31258_ (.A(_08910_),
    .B(_08911_),
    .Y(_08917_));
 sky130_fd_sc_hd__nand3_2 _31259_ (.A(_08916_),
    .B(_08913_),
    .C(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__a21oi_2 _31260_ (.A1(_08547_),
    .A2(_08544_),
    .B1(_08552_),
    .Y(_08919_));
 sky130_fd_sc_hd__nand3_4 _31261_ (.A(_08915_),
    .B(_08918_),
    .C(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__o21ai_2 _31262_ (.A1(_08909_),
    .A2(_08912_),
    .B1(_08913_),
    .Y(_08921_));
 sky130_fd_sc_hd__nand3_2 _31263_ (.A(_08916_),
    .B(_08914_),
    .C(_08917_),
    .Y(_08922_));
 sky130_fd_sc_hd__o21ai_2 _31264_ (.A1(_08546_),
    .A2(_08551_),
    .B1(_08542_),
    .Y(_08923_));
 sky130_fd_sc_hd__nand3_4 _31265_ (.A(_08921_),
    .B(_08922_),
    .C(_08923_),
    .Y(_08924_));
 sky130_fd_sc_hd__a22oi_4 _31266_ (.A1(_19621_),
    .A2(_05268_),
    .B1(_08172_),
    .B2(_05637_),
    .Y(_08925_));
 sky130_fd_sc_hd__nand2_2 _31267_ (.A(_19620_),
    .B(_19916_),
    .Y(_08926_));
 sky130_fd_sc_hd__nand2_2 _31268_ (.A(_07824_),
    .B(_05483_),
    .Y(_08927_));
 sky130_fd_sc_hd__nor2_4 _31269_ (.A(_08926_),
    .B(_08927_),
    .Y(_08928_));
 sky130_fd_sc_hd__nand2_2 _31270_ (.A(_07481_),
    .B(_05769_),
    .Y(_08929_));
 sky130_fd_sc_hd__o21bai_2 _31271_ (.A1(_08925_),
    .A2(_08928_),
    .B1_N(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__nand3b_4 _31272_ (.A_N(_08926_),
    .B(_08567_),
    .C(_05380_),
    .Y(_08931_));
 sky130_fd_sc_hd__nand2_2 _31273_ (.A(_08926_),
    .B(_08927_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand3_2 _31274_ (.A(_08931_),
    .B(_08929_),
    .C(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__nand2_4 _31275_ (.A(_08930_),
    .B(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__nand3_2 _31276_ (.A(_08920_),
    .B(_08924_),
    .C(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__nand2_1 _31277_ (.A(_08920_),
    .B(_08924_),
    .Y(_08936_));
 sky130_vsdinv _31278_ (.A(_08934_),
    .Y(_08937_));
 sky130_fd_sc_hd__nand2_1 _31279_ (.A(_08936_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__nand3_4 _31280_ (.A(_08907_),
    .B(_08935_),
    .C(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__a21boi_4 _31281_ (.A1(_08558_),
    .A2(_08570_),
    .B1_N(_08554_),
    .Y(_08940_));
 sky130_fd_sc_hd__nand2_1 _31282_ (.A(_08936_),
    .B(_08934_),
    .Y(_08941_));
 sky130_fd_sc_hd__nand3_2 _31283_ (.A(_08937_),
    .B(_08920_),
    .C(_08924_),
    .Y(_08942_));
 sky130_fd_sc_hd__nand3_4 _31284_ (.A(_08940_),
    .B(_08941_),
    .C(_08942_),
    .Y(_08943_));
 sky130_fd_sc_hd__nand2_2 _31285_ (.A(_08939_),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__clkbuf_4 _31286_ (.A(\pcpi_mul.rs2[25] ),
    .X(_08945_));
 sky130_fd_sc_hd__clkbuf_4 _31287_ (.A(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__buf_6 _31288_ (.A(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__nand2_1 _31289_ (.A(_08947_),
    .B(_05213_),
    .Y(_08948_));
 sky130_fd_sc_hd__nand2_4 _31290_ (.A(_19603_),
    .B(_05158_),
    .Y(_08949_));
 sky130_fd_sc_hd__nor2_2 _31291_ (.A(_08948_),
    .B(_08949_),
    .Y(_08950_));
 sky130_fd_sc_hd__and2_1 _31292_ (.A(_08948_),
    .B(_08949_),
    .X(_08951_));
 sky130_fd_sc_hd__nor2_4 _31293_ (.A(_08950_),
    .B(_08951_),
    .Y(_08952_));
 sky130_vsdinv _31294_ (.A(_08952_),
    .Y(_08953_));
 sky130_fd_sc_hd__nand2_4 _31295_ (.A(_08944_),
    .B(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__nand3_4 _31296_ (.A(_08939_),
    .B(_08943_),
    .C(_08952_),
    .Y(_08955_));
 sky130_fd_sc_hd__a21boi_1 _31297_ (.A1(_08954_),
    .A2(_08955_),
    .B1_N(_08584_),
    .Y(_08956_));
 sky130_fd_sc_hd__nand2_4 _31298_ (.A(_08954_),
    .B(_08955_),
    .Y(_08957_));
 sky130_fd_sc_hd__nor2_4 _31299_ (.A(_08584_),
    .B(_08957_),
    .Y(_08958_));
 sky130_fd_sc_hd__nor2_2 _31300_ (.A(_08956_),
    .B(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__o21ai_2 _31301_ (.A1(_08904_),
    .A2(_08906_),
    .B1(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__nor2_4 _31302_ (.A(_08636_),
    .B(_08838_),
    .Y(_08961_));
 sky130_fd_sc_hd__a21o_1 _31303_ (.A1(_08903_),
    .A2(_08898_),
    .B1(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__nand3_1 _31304_ (.A(_08663_),
    .B(_08954_),
    .C(_08955_),
    .Y(_08963_));
 sky130_fd_sc_hd__nand2_2 _31305_ (.A(_08957_),
    .B(_08584_),
    .Y(_08964_));
 sky130_fd_sc_hd__nand2_1 _31306_ (.A(_08963_),
    .B(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__nand3_4 _31307_ (.A(_08903_),
    .B(_08898_),
    .C(_08961_),
    .Y(_08966_));
 sky130_fd_sc_hd__nand3_2 _31308_ (.A(_08962_),
    .B(_08965_),
    .C(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__nand3_4 _31309_ (.A(_08960_),
    .B(_08659_),
    .C(_08967_),
    .Y(_08968_));
 sky130_fd_sc_hd__o21ai_2 _31310_ (.A1(_08904_),
    .A2(_08906_),
    .B1(_08965_),
    .Y(_08969_));
 sky130_fd_sc_hd__nand3_2 _31311_ (.A(_08959_),
    .B(_08962_),
    .C(_08966_),
    .Y(_08970_));
 sky130_fd_sc_hd__nand3_4 _31312_ (.A(_08969_),
    .B(_08672_),
    .C(_08970_),
    .Y(_08971_));
 sky130_fd_sc_hd__nand2_1 _31313_ (.A(_08968_),
    .B(_08971_),
    .Y(_08972_));
 sky130_fd_sc_hd__nand2_1 _31314_ (.A(_08837_),
    .B(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__and3_1 _31315_ (.A(_08826_),
    .B(_08828_),
    .C(_08831_),
    .X(_08974_));
 sky130_fd_sc_hd__nand2_4 _31316_ (.A(_08823_),
    .B(_08835_),
    .Y(_08975_));
 sky130_fd_sc_hd__o2111ai_4 _31317_ (.A1(_08974_),
    .A2(_08975_),
    .B1(_08968_),
    .C1(_08971_),
    .D1(_08834_),
    .Y(_08976_));
 sky130_fd_sc_hd__nand3_4 _31318_ (.A(_08729_),
    .B(_08973_),
    .C(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__and3_1 _31319_ (.A(_08383_),
    .B(_08667_),
    .C(_08659_),
    .X(_08978_));
 sky130_fd_sc_hd__a31oi_4 _31320_ (.A1(_08676_),
    .A2(_08673_),
    .A3(_08677_),
    .B1(_08978_),
    .Y(_08979_));
 sky130_fd_sc_hd__nand3_2 _31321_ (.A(_08837_),
    .B(_08968_),
    .C(_08971_),
    .Y(_08980_));
 sky130_fd_sc_hd__nand3_2 _31322_ (.A(_08972_),
    .B(_08834_),
    .C(_08836_),
    .Y(_08981_));
 sky130_fd_sc_hd__nand3_4 _31323_ (.A(_08979_),
    .B(_08980_),
    .C(_08981_),
    .Y(_08982_));
 sky130_fd_sc_hd__nand2_1 _31324_ (.A(_08977_),
    .B(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__a31o_1 _31325_ (.A1(_08499_),
    .A2(_08497_),
    .A3(_08503_),
    .B1(_08509_),
    .X(_08984_));
 sky130_vsdinv _31326_ (.A(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__a21oi_4 _31327_ (.A1(_08684_),
    .A2(_08530_),
    .B1(_08985_),
    .Y(_08986_));
 sky130_fd_sc_hd__and3_2 _31328_ (.A(_08684_),
    .B(_08530_),
    .C(_08985_),
    .X(_08987_));
 sky130_fd_sc_hd__nor2_8 _31329_ (.A(_08986_),
    .B(_08987_),
    .Y(_08988_));
 sky130_fd_sc_hd__nand2_1 _31330_ (.A(_08983_),
    .B(_08988_),
    .Y(_08989_));
 sky130_fd_sc_hd__a21oi_4 _31331_ (.A1(_08670_),
    .A2(_08678_),
    .B1(_08440_),
    .Y(_08990_));
 sky130_fd_sc_hd__a21oi_4 _31332_ (.A1(_08679_),
    .A2(_08697_),
    .B1(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__nand3b_4 _31333_ (.A_N(_08988_),
    .B(_08977_),
    .C(_08982_),
    .Y(_08992_));
 sky130_fd_sc_hd__nand3_4 _31334_ (.A(_08989_),
    .B(_08991_),
    .C(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__a31oi_4 _31335_ (.A1(_08440_),
    .A2(_08670_),
    .A3(_08678_),
    .B1(_08693_),
    .Y(_08994_));
 sky130_fd_sc_hd__nand3_4 _31336_ (.A(_08977_),
    .B(_08982_),
    .C(_08988_),
    .Y(_08995_));
 sky130_fd_sc_hd__o2bb2ai_2 _31337_ (.A1_N(_08982_),
    .A2_N(_08977_),
    .B1(_08986_),
    .B2(_08987_),
    .Y(_08996_));
 sky130_fd_sc_hd__o211ai_4 _31338_ (.A1(_08990_),
    .A2(_08994_),
    .B1(_08995_),
    .C1(_08996_),
    .Y(_08997_));
 sky130_fd_sc_hd__nand2_1 _31339_ (.A(_08993_),
    .B(_08997_),
    .Y(_08998_));
 sky130_vsdinv _31340_ (.A(_08690_),
    .Y(_08999_));
 sky130_fd_sc_hd__nand2_1 _31341_ (.A(_08998_),
    .B(_08999_),
    .Y(_09000_));
 sky130_fd_sc_hd__a21oi_4 _31342_ (.A1(_08679_),
    .A2(_08686_),
    .B1(_08697_),
    .Y(_09001_));
 sky130_fd_sc_hd__and3_1 _31343_ (.A(_08150_),
    .B(_08381_),
    .C(_08388_),
    .X(_09002_));
 sky130_fd_sc_hd__a31oi_2 _31344_ (.A1(_08392_),
    .A2(_08393_),
    .A3(_08394_),
    .B1(_08408_),
    .Y(_09003_));
 sky130_fd_sc_hd__o21ai_2 _31345_ (.A1(_09002_),
    .A2(_09003_),
    .B1(_08698_),
    .Y(_09004_));
 sky130_fd_sc_hd__a2bb2oi_4 _31346_ (.A1_N(_09001_),
    .A2_N(_09004_),
    .B1(_08411_),
    .B2(_08706_),
    .Y(_09005_));
 sky130_fd_sc_hd__nand3_2 _31347_ (.A(_08993_),
    .B(_08997_),
    .C(_08690_),
    .Y(_09006_));
 sky130_fd_sc_hd__nand3_4 _31348_ (.A(_09000_),
    .B(_09005_),
    .C(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__o2bb2ai_1 _31349_ (.A1_N(_08997_),
    .A2_N(_08993_),
    .B1(_08691_),
    .B2(_08700_),
    .Y(_09008_));
 sky130_fd_sc_hd__o2bb2ai_2 _31350_ (.A1_N(_08411_),
    .A2_N(_08706_),
    .B1(_09001_),
    .B2(_09004_),
    .Y(_09009_));
 sky130_fd_sc_hd__nand3_2 _31351_ (.A(_08993_),
    .B(_08997_),
    .C(_08999_),
    .Y(_09010_));
 sky130_fd_sc_hd__nand3_4 _31352_ (.A(_09008_),
    .B(_09009_),
    .C(_09010_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand2_4 _31353_ (.A(_09007_),
    .B(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__o21a_1 _31354_ (.A1(_08717_),
    .A2(_08726_),
    .B1(_08716_),
    .X(_09013_));
 sky130_fd_sc_hd__xor2_4 _31355_ (.A(_09012_),
    .B(_09013_),
    .X(_02644_));
 sky130_fd_sc_hd__nand2_1 _31356_ (.A(_08818_),
    .B(_08805_),
    .Y(_09014_));
 sky130_vsdinv _31357_ (.A(_09014_),
    .Y(_09015_));
 sky130_fd_sc_hd__a21oi_4 _31358_ (.A1(_08975_),
    .A2(_08832_),
    .B1(_09015_),
    .Y(_09016_));
 sky130_fd_sc_hd__and3_2 _31359_ (.A(_08975_),
    .B(_08832_),
    .C(_09015_),
    .X(_09017_));
 sky130_vsdinv _31360_ (.A(_08743_),
    .Y(_09018_));
 sky130_fd_sc_hd__nor2_2 _31361_ (.A(_08750_),
    .B(_08757_),
    .Y(_09019_));
 sky130_fd_sc_hd__a22oi_4 _31362_ (.A1(_05446_),
    .A2(_19873_),
    .B1(_05447_),
    .B2(_07702_),
    .Y(_09020_));
 sky130_fd_sc_hd__and4_4 _31363_ (.A(_05446_),
    .B(_05404_),
    .C(_08061_),
    .D(_19873_),
    .X(_09021_));
 sky130_fd_sc_hd__nand2_2 _31364_ (.A(_05443_),
    .B(_07542_),
    .Y(_09022_));
 sky130_fd_sc_hd__o21ai_2 _31365_ (.A1(_09020_),
    .A2(_09021_),
    .B1(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__nand2_1 _31366_ (.A(_05591_),
    .B(_07345_),
    .Y(_09024_));
 sky130_fd_sc_hd__nand3b_4 _31367_ (.A_N(_09024_),
    .B(_06835_),
    .C(_19871_),
    .Y(_09025_));
 sky130_vsdinv _31368_ (.A(_09022_),
    .Y(_09026_));
 sky130_fd_sc_hd__a22o_1 _31369_ (.A1(_06492_),
    .A2(_19873_),
    .B1(_06217_),
    .B2(_07325_),
    .X(_09027_));
 sky130_fd_sc_hd__nand3_2 _31370_ (.A(_09025_),
    .B(_09026_),
    .C(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__o21ai_2 _31371_ (.A1(_08858_),
    .A2(_08854_),
    .B1(_08860_),
    .Y(_09029_));
 sky130_fd_sc_hd__nand3_4 _31372_ (.A(_09023_),
    .B(_09028_),
    .C(_09029_),
    .Y(_09030_));
 sky130_fd_sc_hd__o21ai_2 _31373_ (.A1(_09020_),
    .A2(_09021_),
    .B1(_09026_),
    .Y(_09031_));
 sky130_fd_sc_hd__nand3_2 _31374_ (.A(_09025_),
    .B(_09022_),
    .C(_09027_),
    .Y(_09032_));
 sky130_fd_sc_hd__o21ai_1 _31375_ (.A1(_08855_),
    .A2(_08856_),
    .B1(_08858_),
    .Y(_09033_));
 sky130_fd_sc_hd__nand2_1 _31376_ (.A(_09033_),
    .B(_08861_),
    .Y(_09034_));
 sky130_fd_sc_hd__nand3_4 _31377_ (.A(_09031_),
    .B(_09032_),
    .C(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__nor2_4 _31378_ (.A(_08741_),
    .B(_08732_),
    .Y(_09036_));
 sky130_fd_sc_hd__o2bb2ai_4 _31379_ (.A1_N(_09030_),
    .A2_N(_09035_),
    .B1(_08740_),
    .B2(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__nor2_4 _31380_ (.A(_08740_),
    .B(_09036_),
    .Y(_09038_));
 sky130_fd_sc_hd__nand3_4 _31381_ (.A(_09030_),
    .B(_09035_),
    .C(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__nand2_1 _31382_ (.A(_08853_),
    .B(_08863_),
    .Y(_09040_));
 sky130_fd_sc_hd__nand2_4 _31383_ (.A(_09040_),
    .B(_08850_),
    .Y(_09041_));
 sky130_fd_sc_hd__a21oi_4 _31384_ (.A1(_09037_),
    .A2(_09039_),
    .B1(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__and3_1 _31385_ (.A(_09041_),
    .B(_09037_),
    .C(_09039_),
    .X(_09043_));
 sky130_fd_sc_hd__o22ai_4 _31386_ (.A1(_09018_),
    .A2(_09019_),
    .B1(_09042_),
    .B2(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__and2_1 _31387_ (.A(_08758_),
    .B(_08748_),
    .X(_09045_));
 sky130_fd_sc_hd__a21o_1 _31388_ (.A1(_09037_),
    .A2(_09039_),
    .B1(_09041_),
    .X(_09046_));
 sky130_fd_sc_hd__nand3_4 _31389_ (.A(_09041_),
    .B(_09037_),
    .C(_09039_),
    .Y(_09047_));
 sky130_fd_sc_hd__nand3b_2 _31390_ (.A_N(_09045_),
    .B(_09046_),
    .C(_09047_),
    .Y(_09048_));
 sky130_vsdinv _31391_ (.A(_08752_),
    .Y(_09049_));
 sky130_fd_sc_hd__nand2_1 _31392_ (.A(_08755_),
    .B(_08751_),
    .Y(_09050_));
 sky130_fd_sc_hd__o22ai_4 _31393_ (.A1(_09049_),
    .A2(_09050_),
    .B1(_08764_),
    .B2(_08756_),
    .Y(_09051_));
 sky130_fd_sc_hd__nand3_4 _31394_ (.A(_09044_),
    .B(_09048_),
    .C(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__o21bai_2 _31395_ (.A1(_09042_),
    .A2(_09043_),
    .B1_N(_09045_),
    .Y(_09053_));
 sky130_fd_sc_hd__nand2_1 _31396_ (.A(_08763_),
    .B(_08764_),
    .Y(_09054_));
 sky130_fd_sc_hd__nand2_1 _31397_ (.A(_09054_),
    .B(_08762_),
    .Y(_09055_));
 sky130_fd_sc_hd__nand3_2 _31398_ (.A(_09046_),
    .B(_09047_),
    .C(_09045_),
    .Y(_09056_));
 sky130_fd_sc_hd__nand3_4 _31399_ (.A(_09053_),
    .B(_09055_),
    .C(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__nand2_2 _31400_ (.A(_05203_),
    .B(_19865_),
    .Y(_09058_));
 sky130_fd_sc_hd__nand2_2 _31401_ (.A(_05366_),
    .B(_08331_),
    .Y(_09059_));
 sky130_fd_sc_hd__nor2_4 _31402_ (.A(_09058_),
    .B(_09059_),
    .Y(_09060_));
 sky130_vsdinv _31403_ (.A(_09060_),
    .Y(_09061_));
 sky130_fd_sc_hd__nand2_4 _31404_ (.A(net495),
    .B(_19847_),
    .Y(_09062_));
 sky130_vsdinv _31405_ (.A(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__nand2_2 _31406_ (.A(_09058_),
    .B(_09059_),
    .Y(_09064_));
 sky130_fd_sc_hd__nand3_2 _31407_ (.A(_09061_),
    .B(_09063_),
    .C(_09064_),
    .Y(_09065_));
 sky130_fd_sc_hd__o21ai_1 _31408_ (.A1(_08782_),
    .A2(_08783_),
    .B1(_08788_),
    .Y(_09066_));
 sky130_fd_sc_hd__and2_1 _31409_ (.A(_09066_),
    .B(_08785_),
    .X(_09067_));
 sky130_fd_sc_hd__a22oi_4 _31410_ (.A1(net455),
    .A2(_19866_),
    .B1(_05780_),
    .B2(_19863_),
    .Y(_09068_));
 sky130_fd_sc_hd__o21ai_2 _31411_ (.A1(_09068_),
    .A2(_09060_),
    .B1(_09062_),
    .Y(_09069_));
 sky130_fd_sc_hd__nand3_4 _31412_ (.A(_09065_),
    .B(_09067_),
    .C(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__nand3_2 _31413_ (.A(_09061_),
    .B(_09062_),
    .C(_09064_),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_1 _31414_ (.A(_09066_),
    .B(_08785_),
    .Y(_09072_));
 sky130_fd_sc_hd__o21ai_2 _31415_ (.A1(_09068_),
    .A2(_09060_),
    .B1(_09063_),
    .Y(_09073_));
 sky130_fd_sc_hd__nand3_4 _31416_ (.A(_09071_),
    .B(_09072_),
    .C(_09073_),
    .Y(_09074_));
 sky130_fd_sc_hd__buf_6 _31417_ (.A(\pcpi_mul.rs1[25] ),
    .X(_09075_));
 sky130_fd_sc_hd__clkbuf_4 _31418_ (.A(\pcpi_mul.rs1[24] ),
    .X(_09076_));
 sky130_fd_sc_hd__nand2_1 _31419_ (.A(_05161_),
    .B(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__a21o_1 _31420_ (.A1(_05239_),
    .A2(_09075_),
    .B1(_09077_),
    .X(_09078_));
 sky130_fd_sc_hd__clkbuf_4 _31421_ (.A(\pcpi_mul.rs1[25] ),
    .X(_09079_));
 sky130_fd_sc_hd__nand2_1 _31422_ (.A(_05382_),
    .B(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__a21o_1 _31423_ (.A1(_06636_),
    .A2(_19854_),
    .B1(_09080_),
    .X(_09081_));
 sky130_fd_sc_hd__buf_6 _31424_ (.A(_08477_),
    .X(_09082_));
 sky130_fd_sc_hd__nand2_2 _31425_ (.A(_05670_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__a21oi_4 _31426_ (.A1(_09078_),
    .A2(_09081_),
    .B1(_09083_),
    .Y(_09084_));
 sky130_fd_sc_hd__and3_2 _31427_ (.A(_09078_),
    .B(_09081_),
    .C(_09083_),
    .X(_09085_));
 sky130_fd_sc_hd__nor2_8 _31428_ (.A(_09084_),
    .B(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__a21o_1 _31429_ (.A1(_09070_),
    .A2(_09074_),
    .B1(_09086_),
    .X(_09087_));
 sky130_fd_sc_hd__nand3_4 _31430_ (.A(_09086_),
    .B(_09070_),
    .C(_09074_),
    .Y(_09088_));
 sky130_fd_sc_hd__nand2_1 _31431_ (.A(_08781_),
    .B(_08794_),
    .Y(_09089_));
 sky130_fd_sc_hd__nand2_2 _31432_ (.A(_09089_),
    .B(_08798_),
    .Y(_09090_));
 sky130_fd_sc_hd__a21o_1 _31433_ (.A1(_09087_),
    .A2(_09088_),
    .B1(_09090_),
    .X(_09091_));
 sky130_fd_sc_hd__nand3_2 _31434_ (.A(_09090_),
    .B(_09087_),
    .C(_09088_),
    .Y(_09092_));
 sky130_vsdinv _31435_ (.A(_08802_),
    .Y(_09093_));
 sky130_fd_sc_hd__or2_2 _31436_ (.A(_08774_),
    .B(_09093_),
    .X(_09094_));
 sky130_fd_sc_hd__a21oi_2 _31437_ (.A1(_09091_),
    .A2(_09092_),
    .B1(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__and3_1 _31438_ (.A(_09090_),
    .B(_09087_),
    .C(_09088_),
    .X(_09096_));
 sky130_fd_sc_hd__nand2_1 _31439_ (.A(_09091_),
    .B(_09094_),
    .Y(_09097_));
 sky130_fd_sc_hd__nor2_2 _31440_ (.A(_09096_),
    .B(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__o2bb2ai_4 _31441_ (.A1_N(_09052_),
    .A2_N(_09057_),
    .B1(_09095_),
    .B2(_09098_),
    .Y(_09099_));
 sky130_fd_sc_hd__a21oi_1 _31442_ (.A1(_09087_),
    .A2(_09088_),
    .B1(_09090_),
    .Y(_09100_));
 sky130_fd_sc_hd__o22ai_2 _31443_ (.A1(_08774_),
    .A2(_09093_),
    .B1(_09100_),
    .B2(_09096_),
    .Y(_09101_));
 sky130_fd_sc_hd__nand3b_1 _31444_ (.A_N(_09094_),
    .B(_09091_),
    .C(_09092_),
    .Y(_09102_));
 sky130_fd_sc_hd__nand2_2 _31445_ (.A(_09101_),
    .B(_09102_),
    .Y(_09103_));
 sky130_fd_sc_hd__nand3_4 _31446_ (.A(_09103_),
    .B(_09052_),
    .C(_09057_),
    .Y(_09104_));
 sky130_fd_sc_hd__nand2_2 _31447_ (.A(_09099_),
    .B(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__nor2_2 _31448_ (.A(_08639_),
    .B(_08905_),
    .Y(_09106_));
 sky130_fd_sc_hd__a31oi_4 _31449_ (.A1(_08899_),
    .A2(_08902_),
    .A3(_08573_),
    .B1(_09106_),
    .Y(_09107_));
 sky130_vsdinv _31450_ (.A(_08898_),
    .Y(_09108_));
 sky130_fd_sc_hd__nor2_2 _31451_ (.A(_09107_),
    .B(_09108_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand2_1 _31452_ (.A(_09105_),
    .B(_09109_),
    .Y(_09110_));
 sky130_fd_sc_hd__nand2_1 _31453_ (.A(_08903_),
    .B(_08961_),
    .Y(_09111_));
 sky130_fd_sc_hd__nand2_2 _31454_ (.A(_09111_),
    .B(_08898_),
    .Y(_09112_));
 sky130_fd_sc_hd__nand3_4 _31455_ (.A(_09112_),
    .B(_09099_),
    .C(_09104_),
    .Y(_09113_));
 sky130_vsdinv _31456_ (.A(_08770_),
    .Y(_09114_));
 sky130_fd_sc_hd__a21o_1 _31457_ (.A1(_08766_),
    .A2(_08830_),
    .B1(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__nand3_4 _31458_ (.A(_09110_),
    .B(_09113_),
    .C(_09115_),
    .Y(_09116_));
 sky130_fd_sc_hd__a21oi_2 _31459_ (.A1(_09099_),
    .A2(_09104_),
    .B1(_09112_),
    .Y(_09117_));
 sky130_fd_sc_hd__o211a_2 _31460_ (.A1(_09107_),
    .A2(_09108_),
    .B1(_09104_),
    .C1(_09099_),
    .X(_09118_));
 sky130_fd_sc_hd__o21bai_4 _31461_ (.A1(_09117_),
    .A2(_09118_),
    .B1_N(_09115_),
    .Y(_09119_));
 sky130_fd_sc_hd__nand2_2 _31462_ (.A(_08881_),
    .B(_08882_),
    .Y(_09120_));
 sky130_fd_sc_hd__a22oi_4 _31463_ (.A1(_19631_),
    .A2(_06264_),
    .B1(_19635_),
    .B2(_05798_),
    .Y(_09121_));
 sky130_fd_sc_hd__nand3_4 _31464_ (.A(_07743_),
    .B(_19634_),
    .C(_05801_),
    .Y(_09122_));
 sky130_fd_sc_hd__nor2_8 _31465_ (.A(net446),
    .B(_09122_),
    .Y(_09123_));
 sky130_fd_sc_hd__nand2_2 _31466_ (.A(_19640_),
    .B(_19897_),
    .Y(_09124_));
 sky130_vsdinv _31467_ (.A(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__o21ai_4 _31468_ (.A1(_09121_),
    .A2(_09123_),
    .B1(_09125_),
    .Y(_09126_));
 sky130_vsdinv _31469_ (.A(_08929_),
    .Y(_09127_));
 sky130_fd_sc_hd__a21oi_4 _31470_ (.A1(_09127_),
    .A2(_08932_),
    .B1(_08928_),
    .Y(_09128_));
 sky130_fd_sc_hd__a22o_2 _31471_ (.A1(_06986_),
    .A2(_06826_),
    .B1(_07428_),
    .B2(_06448_),
    .X(_09129_));
 sky130_fd_sc_hd__o211ai_4 _31472_ (.A1(net446),
    .A2(_09122_),
    .B1(_09124_),
    .C1(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__nand3_4 _31473_ (.A(_09126_),
    .B(_09128_),
    .C(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__o21ai_2 _31474_ (.A1(_09121_),
    .A2(_09123_),
    .B1(_09124_),
    .Y(_09132_));
 sky130_fd_sc_hd__o21ai_2 _31475_ (.A1(_08929_),
    .A2(_08925_),
    .B1(_08931_),
    .Y(_09133_));
 sky130_fd_sc_hd__o211ai_2 _31476_ (.A1(net442),
    .A2(_09122_),
    .B1(_09125_),
    .C1(_09129_),
    .Y(_09134_));
 sky130_fd_sc_hd__nand3_4 _31477_ (.A(_09132_),
    .B(_09133_),
    .C(_09134_),
    .Y(_09135_));
 sky130_fd_sc_hd__nor2_2 _31478_ (.A(_08875_),
    .B(_08868_),
    .Y(_09136_));
 sky130_fd_sc_hd__o2bb2ai_4 _31479_ (.A1_N(_09131_),
    .A2_N(_09135_),
    .B1(_08874_),
    .B2(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__o21ai_4 _31480_ (.A1(_08875_),
    .A2(_08868_),
    .B1(_08870_),
    .Y(_09138_));
 sky130_vsdinv _31481_ (.A(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__nand3_4 _31482_ (.A(_09139_),
    .B(_09131_),
    .C(_09135_),
    .Y(_09140_));
 sky130_fd_sc_hd__a22oi_4 _31483_ (.A1(_08877_),
    .A2(_09120_),
    .B1(_09137_),
    .B2(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__a21oi_4 _31484_ (.A1(_09131_),
    .A2(_09135_),
    .B1(_09139_),
    .Y(_09142_));
 sky130_fd_sc_hd__nand3_4 _31485_ (.A(_09140_),
    .B(_08877_),
    .C(_09120_),
    .Y(_09143_));
 sky130_fd_sc_hd__nor2_8 _31486_ (.A(_09142_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__a21oi_4 _31487_ (.A1(_08848_),
    .A2(_08847_),
    .B1(_08842_),
    .Y(_09145_));
 sky130_fd_sc_hd__a22oi_4 _31488_ (.A1(_06341_),
    .A2(_06788_),
    .B1(_06422_),
    .B2(_07281_),
    .Y(_09146_));
 sky130_fd_sc_hd__nand2_2 _31489_ (.A(_06605_),
    .B(_06115_),
    .Y(_09147_));
 sky130_fd_sc_hd__nand2_2 _31490_ (.A(_06168_),
    .B(_06779_),
    .Y(_09148_));
 sky130_fd_sc_hd__nor2_4 _31491_ (.A(_09147_),
    .B(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__nand2_2 _31492_ (.A(_07223_),
    .B(_19887_),
    .Y(_09150_));
 sky130_vsdinv _31493_ (.A(_09150_),
    .Y(_09151_));
 sky130_fd_sc_hd__o21ai_2 _31494_ (.A1(_09146_),
    .A2(_09149_),
    .B1(_09151_),
    .Y(_09152_));
 sky130_fd_sc_hd__nand3b_4 _31495_ (.A_N(_09147_),
    .B(_06898_),
    .C(_06780_),
    .Y(_09153_));
 sky130_fd_sc_hd__nand2_2 _31496_ (.A(_09147_),
    .B(_09148_),
    .Y(_09154_));
 sky130_fd_sc_hd__nand3_2 _31497_ (.A(_09153_),
    .B(_09150_),
    .C(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__nand3_4 _31498_ (.A(_09145_),
    .B(_09152_),
    .C(_09155_),
    .Y(_09156_));
 sky130_vsdinv _31499_ (.A(_09156_),
    .Y(_09157_));
 sky130_fd_sc_hd__o21ai_2 _31500_ (.A1(_09146_),
    .A2(_09149_),
    .B1(_09150_),
    .Y(_09158_));
 sky130_fd_sc_hd__nand3_2 _31501_ (.A(_09153_),
    .B(_09151_),
    .C(_09154_),
    .Y(_09159_));
 sky130_fd_sc_hd__o21ai_2 _31502_ (.A1(_08843_),
    .A2(_08841_),
    .B1(_08846_),
    .Y(_09160_));
 sky130_fd_sc_hd__nand3_4 _31503_ (.A(_09158_),
    .B(_09159_),
    .C(_09160_),
    .Y(_09161_));
 sky130_fd_sc_hd__a22oi_4 _31504_ (.A1(_07893_),
    .A2(_07059_),
    .B1(_06884_),
    .B2(_08280_),
    .Y(_09162_));
 sky130_fd_sc_hd__nand2_2 _31505_ (.A(_06882_),
    .B(_19883_),
    .Y(_09163_));
 sky130_fd_sc_hd__nand2_1 _31506_ (.A(_06024_),
    .B(_06803_),
    .Y(_09164_));
 sky130_fd_sc_hd__nor2_2 _31507_ (.A(_09163_),
    .B(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__nand2_2 _31508_ (.A(_05731_),
    .B(_06783_),
    .Y(_09166_));
 sky130_fd_sc_hd__o21bai_1 _31509_ (.A1(_09162_),
    .A2(_09165_),
    .B1_N(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__nand3b_4 _31510_ (.A_N(_09163_),
    .B(_06159_),
    .C(_19881_),
    .Y(_09168_));
 sky130_fd_sc_hd__nand2_1 _31511_ (.A(_09163_),
    .B(_09164_),
    .Y(_09169_));
 sky130_fd_sc_hd__nand3_2 _31512_ (.A(_09168_),
    .B(_09166_),
    .C(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__nand2_1 _31513_ (.A(_09167_),
    .B(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__nand2_2 _31514_ (.A(_09161_),
    .B(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__a21o_1 _31515_ (.A1(_09156_),
    .A2(_09161_),
    .B1(_09171_),
    .X(_09173_));
 sky130_fd_sc_hd__o21ai_4 _31516_ (.A1(_09157_),
    .A2(_09172_),
    .B1(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__o21ai_2 _31517_ (.A1(_09141_),
    .A2(_09144_),
    .B1(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__nand2_1 _31518_ (.A(_08890_),
    .B(_08881_),
    .Y(_09176_));
 sky130_fd_sc_hd__a21o_1 _31519_ (.A1(_09137_),
    .A2(_09140_),
    .B1(_09176_),
    .X(_09177_));
 sky130_fd_sc_hd__nand3_2 _31520_ (.A(_09176_),
    .B(_09137_),
    .C(_09140_),
    .Y(_09178_));
 sky130_fd_sc_hd__o21a_2 _31521_ (.A1(_09157_),
    .A2(_09172_),
    .B1(_09173_),
    .X(_09179_));
 sky130_fd_sc_hd__nand3_2 _31522_ (.A(_09177_),
    .B(_09178_),
    .C(_09179_),
    .Y(_09180_));
 sky130_vsdinv _31523_ (.A(_08939_),
    .Y(_09181_));
 sky130_fd_sc_hd__nand3_4 _31524_ (.A(_09175_),
    .B(_09180_),
    .C(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__o21ai_2 _31525_ (.A1(_09141_),
    .A2(_09144_),
    .B1(_09179_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand3_2 _31526_ (.A(_09177_),
    .B(_09178_),
    .C(_09174_),
    .Y(_09184_));
 sky130_fd_sc_hd__nand3_4 _31527_ (.A(_09183_),
    .B(_09184_),
    .C(_08939_),
    .Y(_09185_));
 sky130_fd_sc_hd__nand2_1 _31528_ (.A(_08901_),
    .B(_08895_),
    .Y(_09186_));
 sky130_vsdinv _31529_ (.A(_09186_),
    .Y(_09187_));
 sky130_fd_sc_hd__o2bb2ai_4 _31530_ (.A1_N(_09182_),
    .A2_N(_09185_),
    .B1(_08888_),
    .B2(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__and2_2 _31531_ (.A(_09186_),
    .B(_08894_),
    .X(_09189_));
 sky130_fd_sc_hd__nand3_4 _31532_ (.A(_09182_),
    .B(_09185_),
    .C(_09189_),
    .Y(_09190_));
 sky130_fd_sc_hd__buf_4 _31533_ (.A(\pcpi_mul.rs2[23] ),
    .X(_09191_));
 sky130_fd_sc_hd__a22oi_4 _31534_ (.A1(_09191_),
    .A2(_19923_),
    .B1(_08154_),
    .B2(_05272_),
    .Y(_09192_));
 sky130_fd_sc_hd__nand2_2 _31535_ (.A(_19606_),
    .B(_19922_),
    .Y(_09193_));
 sky130_fd_sc_hd__nand2_2 _31536_ (.A(_19610_),
    .B(_19919_),
    .Y(_09194_));
 sky130_fd_sc_hd__nor2_4 _31537_ (.A(_09193_),
    .B(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__nand2_2 _31538_ (.A(_19615_),
    .B(_05267_),
    .Y(_09196_));
 sky130_fd_sc_hd__o21ai_2 _31539_ (.A1(_09192_),
    .A2(_09195_),
    .B1(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__nand3b_4 _31540_ (.A_N(_09193_),
    .B(_19611_),
    .C(_07008_),
    .Y(_09198_));
 sky130_vsdinv _31541_ (.A(_09196_),
    .Y(_09199_));
 sky130_fd_sc_hd__nand2_2 _31542_ (.A(_09193_),
    .B(_09194_),
    .Y(_09200_));
 sky130_fd_sc_hd__nand3_2 _31543_ (.A(_09198_),
    .B(_09199_),
    .C(_09200_),
    .Y(_09201_));
 sky130_fd_sc_hd__o21ai_2 _31544_ (.A1(_08913_),
    .A2(_08909_),
    .B1(_08916_),
    .Y(_09202_));
 sky130_fd_sc_hd__nand3_4 _31545_ (.A(_09197_),
    .B(_09201_),
    .C(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__o21ai_2 _31546_ (.A1(_09192_),
    .A2(_09195_),
    .B1(_09199_),
    .Y(_09204_));
 sky130_fd_sc_hd__nand3_2 _31547_ (.A(_09198_),
    .B(_09196_),
    .C(_09200_),
    .Y(_09205_));
 sky130_fd_sc_hd__a21oi_4 _31548_ (.A1(_08914_),
    .A2(_08917_),
    .B1(_08912_),
    .Y(_09206_));
 sky130_fd_sc_hd__nand3_4 _31549_ (.A(_09204_),
    .B(_09205_),
    .C(_09206_),
    .Y(_09207_));
 sky130_fd_sc_hd__a22oi_4 _31550_ (.A1(_07933_),
    .A2(_05379_),
    .B1(_07258_),
    .B2(_05488_),
    .Y(_09208_));
 sky130_fd_sc_hd__nand2_2 _31551_ (.A(\pcpi_mul.rs2[20] ),
    .B(_19912_),
    .Y(_09209_));
 sky130_fd_sc_hd__nand2_2 _31552_ (.A(_19624_),
    .B(_05480_),
    .Y(_09210_));
 sky130_fd_sc_hd__nor2_4 _31553_ (.A(_09209_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__nand2_2 _31554_ (.A(\pcpi_mul.rs2[18] ),
    .B(_05463_),
    .Y(_09212_));
 sky130_fd_sc_hd__o21a_1 _31555_ (.A1(_09208_),
    .A2(_09211_),
    .B1(_09212_),
    .X(_09213_));
 sky130_fd_sc_hd__nand3b_4 _31556_ (.A_N(_09209_),
    .B(_07827_),
    .C(_05545_),
    .Y(_09214_));
 sky130_vsdinv _31557_ (.A(_09212_),
    .Y(_09215_));
 sky130_fd_sc_hd__nand2_2 _31558_ (.A(_09209_),
    .B(_09210_),
    .Y(_09216_));
 sky130_fd_sc_hd__and3_1 _31559_ (.A(_09214_),
    .B(_09215_),
    .C(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__o2bb2ai_4 _31560_ (.A1_N(_09203_),
    .A2_N(_09207_),
    .B1(_09213_),
    .B2(_09217_),
    .Y(_09218_));
 sky130_fd_sc_hd__o21ai_2 _31561_ (.A1(_09208_),
    .A2(_09211_),
    .B1(_09215_),
    .Y(_09219_));
 sky130_fd_sc_hd__nand3_2 _31562_ (.A(_09214_),
    .B(_09212_),
    .C(_09216_),
    .Y(_09220_));
 sky130_fd_sc_hd__nand2_4 _31563_ (.A(_09219_),
    .B(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__nand3_4 _31564_ (.A(_09207_),
    .B(_09203_),
    .C(_09221_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand2_1 _31565_ (.A(_08920_),
    .B(_08934_),
    .Y(_09223_));
 sky130_fd_sc_hd__nand2_4 _31566_ (.A(_09223_),
    .B(_08924_),
    .Y(_09224_));
 sky130_fd_sc_hd__a21o_1 _31567_ (.A1(_09218_),
    .A2(_09222_),
    .B1(_09224_),
    .X(_09225_));
 sky130_vsdinv _31568_ (.A(_08950_),
    .Y(_09226_));
 sky130_fd_sc_hd__buf_4 _31569_ (.A(_08945_),
    .X(_09227_));
 sky130_fd_sc_hd__nand2_2 _31570_ (.A(_09227_),
    .B(_05122_),
    .Y(_09228_));
 sky130_fd_sc_hd__clkbuf_4 _31571_ (.A(\pcpi_mul.rs2[26] ),
    .X(_09229_));
 sky130_fd_sc_hd__nand2_2 _31572_ (.A(_09229_),
    .B(_19932_),
    .Y(_09230_));
 sky130_fd_sc_hd__nor2_4 _31573_ (.A(_09228_),
    .B(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__and2_1 _31574_ (.A(_09228_),
    .B(_09230_),
    .X(_09232_));
 sky130_fd_sc_hd__nor2_4 _31575_ (.A(_08578_),
    .B(_05150_),
    .Y(_09233_));
 sky130_fd_sc_hd__o21bai_4 _31576_ (.A1(_09231_),
    .A2(_09232_),
    .B1_N(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__nand2_2 _31577_ (.A(_09228_),
    .B(_09230_),
    .Y(_09235_));
 sky130_fd_sc_hd__nand3b_4 _31578_ (.A_N(_09231_),
    .B(_09235_),
    .C(_09233_),
    .Y(_09236_));
 sky130_fd_sc_hd__nand2_8 _31579_ (.A(_09234_),
    .B(_09236_),
    .Y(_09237_));
 sky130_fd_sc_hd__nor2_8 _31580_ (.A(_09226_),
    .B(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__and2_1 _31581_ (.A(_09237_),
    .B(_09226_),
    .X(_09239_));
 sky130_fd_sc_hd__nor2_4 _31582_ (.A(_09238_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__nand3_4 _31583_ (.A(_09224_),
    .B(_09218_),
    .C(_09222_),
    .Y(_09241_));
 sky130_fd_sc_hd__nand3_4 _31584_ (.A(_09225_),
    .B(_09240_),
    .C(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__nand2_1 _31585_ (.A(_09225_),
    .B(_09241_),
    .Y(_09243_));
 sky130_vsdinv _31586_ (.A(_09240_),
    .Y(_09244_));
 sky130_fd_sc_hd__a21oi_4 _31587_ (.A1(_09243_),
    .A2(_09244_),
    .B1(_08955_),
    .Y(_09245_));
 sky130_fd_sc_hd__a21oi_1 _31588_ (.A1(_09218_),
    .A2(_09222_),
    .B1(_09224_),
    .Y(_09246_));
 sky130_fd_sc_hd__nand2_2 _31589_ (.A(_09207_),
    .B(_09221_),
    .Y(_09247_));
 sky130_vsdinv _31590_ (.A(_09203_),
    .Y(_09248_));
 sky130_fd_sc_hd__o211a_1 _31591_ (.A1(_09247_),
    .A2(_09248_),
    .B1(_09218_),
    .C1(_09224_),
    .X(_09249_));
 sky130_fd_sc_hd__o21ai_1 _31592_ (.A1(_09246_),
    .A2(_09249_),
    .B1(_09244_),
    .Y(_09250_));
 sky130_fd_sc_hd__nor2_1 _31593_ (.A(_08953_),
    .B(_08944_),
    .Y(_09251_));
 sky130_fd_sc_hd__a21oi_2 _31594_ (.A1(_09250_),
    .A2(_09242_),
    .B1(_09251_),
    .Y(_09252_));
 sky130_fd_sc_hd__a21oi_4 _31595_ (.A1(_09242_),
    .A2(_09245_),
    .B1(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__a21o_1 _31596_ (.A1(_09188_),
    .A2(_09190_),
    .B1(_09253_),
    .X(_09254_));
 sky130_fd_sc_hd__nand3_4 _31597_ (.A(_09253_),
    .B(_09188_),
    .C(_09190_),
    .Y(_09255_));
 sky130_fd_sc_hd__nand2_1 _31598_ (.A(_08966_),
    .B(_08964_),
    .Y(_09256_));
 sky130_fd_sc_hd__o22ai_4 _31599_ (.A1(_08584_),
    .A2(_08957_),
    .B1(_08904_),
    .B2(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__a21oi_2 _31600_ (.A1(_09254_),
    .A2(_09255_),
    .B1(_09257_),
    .Y(_09258_));
 sky130_vsdinv _31601_ (.A(_09190_),
    .Y(_09259_));
 sky130_fd_sc_hd__nand2_1 _31602_ (.A(_09253_),
    .B(_09188_),
    .Y(_09260_));
 sky130_fd_sc_hd__o211a_2 _31603_ (.A1(_09259_),
    .A2(_09260_),
    .B1(_09254_),
    .C1(_09257_),
    .X(_09261_));
 sky130_fd_sc_hd__o2bb2ai_4 _31604_ (.A1_N(_09116_),
    .A2_N(_09119_),
    .B1(_09258_),
    .B2(_09261_),
    .Y(_09262_));
 sky130_fd_sc_hd__and2_1 _31605_ (.A(_08830_),
    .B(_08766_),
    .X(_09263_));
 sky130_fd_sc_hd__o2bb2ai_4 _31606_ (.A1_N(_09109_),
    .A2_N(_09105_),
    .B1(_09114_),
    .B2(_09263_),
    .Y(_09264_));
 sky130_fd_sc_hd__a21oi_2 _31607_ (.A1(_09188_),
    .A2(_09190_),
    .B1(_09253_),
    .Y(_09265_));
 sky130_vsdinv _31608_ (.A(_09182_),
    .Y(_09266_));
 sky130_fd_sc_hd__nand2_1 _31609_ (.A(_09185_),
    .B(_09189_),
    .Y(_09267_));
 sky130_fd_sc_hd__o211a_1 _31610_ (.A1(_09266_),
    .A2(_09267_),
    .B1(_09188_),
    .C1(_09253_),
    .X(_09268_));
 sky130_fd_sc_hd__a31oi_4 _31611_ (.A1(_08962_),
    .A2(_08966_),
    .A3(_08964_),
    .B1(_08958_),
    .Y(_09269_));
 sky130_fd_sc_hd__o21ai_4 _31612_ (.A1(_09265_),
    .A2(_09268_),
    .B1(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__nand3_4 _31613_ (.A(_09257_),
    .B(_09254_),
    .C(_09255_),
    .Y(_09271_));
 sky130_fd_sc_hd__o2111ai_4 _31614_ (.A1(_09118_),
    .A2(_09264_),
    .B1(_09270_),
    .C1(_09271_),
    .D1(_09119_),
    .Y(_09272_));
 sky130_fd_sc_hd__nand3_2 _31615_ (.A(_08834_),
    .B(_08968_),
    .C(_08836_),
    .Y(_09273_));
 sky130_fd_sc_hd__nand2_4 _31616_ (.A(_09273_),
    .B(_08971_),
    .Y(_09274_));
 sky130_fd_sc_hd__a21oi_4 _31617_ (.A1(_09262_),
    .A2(_09272_),
    .B1(_09274_),
    .Y(_09275_));
 sky130_vsdinv _31618_ (.A(_08971_),
    .Y(_09276_));
 sky130_fd_sc_hd__o211a_1 _31619_ (.A1(_08974_),
    .A2(_08975_),
    .B1(_08968_),
    .C1(_08834_),
    .X(_09277_));
 sky130_fd_sc_hd__o211a_2 _31620_ (.A1(_09276_),
    .A2(_09277_),
    .B1(_09262_),
    .C1(_09272_),
    .X(_09278_));
 sky130_fd_sc_hd__o22ai_4 _31621_ (.A1(_09016_),
    .A2(_09017_),
    .B1(_09275_),
    .B2(_09278_),
    .Y(_09279_));
 sky130_fd_sc_hd__nand2_2 _31622_ (.A(_08995_),
    .B(_08977_),
    .Y(_09280_));
 sky130_fd_sc_hd__a21o_2 _31623_ (.A1(_09262_),
    .A2(_09272_),
    .B1(_09274_),
    .X(_09281_));
 sky130_fd_sc_hd__nand3_4 _31624_ (.A(_09262_),
    .B(_09274_),
    .C(_09272_),
    .Y(_09282_));
 sky130_fd_sc_hd__nor2_8 _31625_ (.A(_09016_),
    .B(_09017_),
    .Y(_09283_));
 sky130_fd_sc_hd__nand3_4 _31626_ (.A(_09281_),
    .B(_09282_),
    .C(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__nand3_4 _31627_ (.A(_09279_),
    .B(_09280_),
    .C(_09284_),
    .Y(_09285_));
 sky130_fd_sc_hd__o21ai_2 _31628_ (.A1(_09275_),
    .A2(_09278_),
    .B1(_09283_),
    .Y(_09286_));
 sky130_fd_sc_hd__a21boi_4 _31629_ (.A1(_08982_),
    .A2(_08988_),
    .B1_N(_08977_),
    .Y(_09287_));
 sky130_vsdinv _31630_ (.A(_09283_),
    .Y(_09288_));
 sky130_fd_sc_hd__nand3_4 _31631_ (.A(_09281_),
    .B(_09282_),
    .C(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__nand3_4 _31632_ (.A(_09286_),
    .B(_09287_),
    .C(_09289_),
    .Y(_09290_));
 sky130_fd_sc_hd__nor2_2 _31633_ (.A(_08683_),
    .B(_08535_),
    .Y(_09291_));
 sky130_fd_sc_hd__o2bb2ai_2 _31634_ (.A1_N(_09285_),
    .A2_N(_09290_),
    .B1(_08985_),
    .B2(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__nand3_2 _31635_ (.A(_09290_),
    .B(_09285_),
    .C(_08986_),
    .Y(_09293_));
 sky130_fd_sc_hd__nand2_1 _31636_ (.A(_08993_),
    .B(_08999_),
    .Y(_09294_));
 sky130_fd_sc_hd__nand2_2 _31637_ (.A(_09294_),
    .B(_08997_),
    .Y(_09295_));
 sky130_fd_sc_hd__a21oi_4 _31638_ (.A1(_09292_),
    .A2(_09293_),
    .B1(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__and3_1 _31639_ (.A(_09279_),
    .B(_09280_),
    .C(_09284_),
    .X(_09297_));
 sky130_fd_sc_hd__nand2_1 _31640_ (.A(_09290_),
    .B(_08986_),
    .Y(_09298_));
 sky130_fd_sc_hd__o211a_2 _31641_ (.A1(_09297_),
    .A2(_09298_),
    .B1(_09295_),
    .C1(_09292_),
    .X(_09299_));
 sky130_fd_sc_hd__nor2_8 _31642_ (.A(_09296_),
    .B(_09299_),
    .Y(_09300_));
 sky130_fd_sc_hd__nand2_4 _31643_ (.A(_08439_),
    .B(_08724_),
    .Y(_09301_));
 sky130_fd_sc_hd__nor2_8 _31644_ (.A(_09012_),
    .B(_08717_),
    .Y(_09302_));
 sky130_fd_sc_hd__a21boi_4 _31645_ (.A1(_08716_),
    .A2(_09011_),
    .B1_N(_09007_),
    .Y(_09303_));
 sky130_fd_sc_hd__a21oi_4 _31646_ (.A1(_09301_),
    .A2(_09302_),
    .B1(_09303_),
    .Y(_09304_));
 sky130_fd_sc_hd__xnor2_2 _31647_ (.A(_09300_),
    .B(_09304_),
    .Y(_02645_));
 sky130_fd_sc_hd__nand3_1 _31648_ (.A(_09119_),
    .B(_09270_),
    .C(_09116_),
    .Y(_09305_));
 sky130_fd_sc_hd__nand2_1 _31649_ (.A(_09305_),
    .B(_09271_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand2_1 _31650_ (.A(_09156_),
    .B(_09171_),
    .Y(_09307_));
 sky130_fd_sc_hd__nand2_2 _31651_ (.A(_09307_),
    .B(_09161_),
    .Y(_09308_));
 sky130_fd_sc_hd__a22oi_4 _31652_ (.A1(_05446_),
    .A2(_07702_),
    .B1(_05447_),
    .B2(_08485_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand3_4 _31653_ (.A(_19661_),
    .B(_05588_),
    .C(_08061_),
    .Y(_09310_));
 sky130_fd_sc_hd__nor2_4 _31654_ (.A(_08078_),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__nand2_2 _31655_ (.A(_05259_),
    .B(_07686_),
    .Y(_09312_));
 sky130_fd_sc_hd__o21ai_2 _31656_ (.A1(_09309_),
    .A2(_09311_),
    .B1(_09312_),
    .Y(_09313_));
 sky130_vsdinv _31657_ (.A(_09312_),
    .Y(_09314_));
 sky130_fd_sc_hd__a22o_1 _31658_ (.A1(_06492_),
    .A2(_07325_),
    .B1(_06217_),
    .B2(_08485_),
    .X(_09315_));
 sky130_fd_sc_hd__o211ai_2 _31659_ (.A1(_08079_),
    .A2(_09310_),
    .B1(_09314_),
    .C1(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__o21ai_2 _31660_ (.A1(_09166_),
    .A2(_09162_),
    .B1(_09168_),
    .Y(_09317_));
 sky130_fd_sc_hd__nand3_4 _31661_ (.A(_09313_),
    .B(_09316_),
    .C(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__o21ai_2 _31662_ (.A1(_09309_),
    .A2(_09311_),
    .B1(_09314_),
    .Y(_09319_));
 sky130_vsdinv _31663_ (.A(_09166_),
    .Y(_09320_));
 sky130_fd_sc_hd__a21oi_2 _31664_ (.A1(_09320_),
    .A2(_09169_),
    .B1(_09165_),
    .Y(_09321_));
 sky130_fd_sc_hd__o211ai_2 _31665_ (.A1(_08079_),
    .A2(_09310_),
    .B1(_09312_),
    .C1(_09315_),
    .Y(_09322_));
 sky130_fd_sc_hd__nand3_4 _31666_ (.A(_09319_),
    .B(_09321_),
    .C(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__nor2_2 _31667_ (.A(_09026_),
    .B(_09021_),
    .Y(_09324_));
 sky130_fd_sc_hd__o2bb2ai_4 _31668_ (.A1_N(_09318_),
    .A2_N(_09323_),
    .B1(_09020_),
    .B2(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__nor2_2 _31669_ (.A(_09022_),
    .B(_09020_),
    .Y(_09326_));
 sky130_fd_sc_hd__o211ai_4 _31670_ (.A1(_09021_),
    .A2(_09326_),
    .B1(_09318_),
    .C1(_09323_),
    .Y(_09327_));
 sky130_fd_sc_hd__nand3_4 _31671_ (.A(_09308_),
    .B(_09325_),
    .C(_09327_),
    .Y(_09328_));
 sky130_fd_sc_hd__and3_1 _31672_ (.A(_09161_),
    .B(_09167_),
    .C(_09170_),
    .X(_09329_));
 sky130_fd_sc_hd__o2bb2ai_4 _31673_ (.A1_N(_09327_),
    .A2_N(_09325_),
    .B1(_09157_),
    .B2(_09329_),
    .Y(_09330_));
 sky130_vsdinv _31674_ (.A(_09030_),
    .Y(_09331_));
 sky130_fd_sc_hd__and2_1 _31675_ (.A(_09035_),
    .B(_09038_),
    .X(_09332_));
 sky130_fd_sc_hd__o2bb2ai_1 _31676_ (.A1_N(_09328_),
    .A2_N(_09330_),
    .B1(_09331_),
    .B2(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__nand2_1 _31677_ (.A(_09047_),
    .B(_09045_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_1 _31678_ (.A(_09334_),
    .B(_09046_),
    .Y(_09335_));
 sky130_fd_sc_hd__nor2_4 _31679_ (.A(_09331_),
    .B(_09332_),
    .Y(_09336_));
 sky130_fd_sc_hd__nand3_2 _31680_ (.A(_09330_),
    .B(_09328_),
    .C(_09336_),
    .Y(_09337_));
 sky130_fd_sc_hd__nand3_4 _31681_ (.A(_09333_),
    .B(_09335_),
    .C(_09337_),
    .Y(_09338_));
 sky130_vsdinv _31682_ (.A(_09035_),
    .Y(_09339_));
 sky130_fd_sc_hd__nor2_1 _31683_ (.A(_09038_),
    .B(_09331_),
    .Y(_09340_));
 sky130_fd_sc_hd__o2bb2ai_1 _31684_ (.A1_N(_09328_),
    .A2_N(_09330_),
    .B1(_09339_),
    .B2(_09340_),
    .Y(_09341_));
 sky130_fd_sc_hd__o21ai_2 _31685_ (.A1(_09045_),
    .A2(_09042_),
    .B1(_09047_),
    .Y(_09342_));
 sky130_fd_sc_hd__nand3b_2 _31686_ (.A_N(_09336_),
    .B(_09330_),
    .C(_09328_),
    .Y(_09343_));
 sky130_fd_sc_hd__nand3_4 _31687_ (.A(_09341_),
    .B(_09342_),
    .C(_09343_),
    .Y(_09344_));
 sky130_fd_sc_hd__nand2_1 _31688_ (.A(_09338_),
    .B(_09344_),
    .Y(_09345_));
 sky130_fd_sc_hd__nand2_2 _31689_ (.A(_19670_),
    .B(_19862_),
    .Y(_09346_));
 sky130_fd_sc_hd__nand2_2 _31690_ (.A(_05282_),
    .B(_08477_),
    .Y(_09347_));
 sky130_fd_sc_hd__or2_4 _31691_ (.A(_09346_),
    .B(_09347_),
    .X(_09348_));
 sky130_fd_sc_hd__a22oi_4 _31692_ (.A1(_05203_),
    .A2(_08331_),
    .B1(_05358_),
    .B2(_08477_),
    .Y(_09349_));
 sky130_vsdinv _31693_ (.A(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__nand2_4 _31694_ (.A(_05290_),
    .B(_19843_),
    .Y(_09351_));
 sky130_vsdinv _31695_ (.A(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand3_4 _31696_ (.A(_09348_),
    .B(_09350_),
    .C(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__nor2_4 _31697_ (.A(_09346_),
    .B(_09347_),
    .Y(_09354_));
 sky130_fd_sc_hd__o21ai_4 _31698_ (.A1(_09349_),
    .A2(_09354_),
    .B1(_09351_),
    .Y(_09355_));
 sky130_fd_sc_hd__a21o_1 _31699_ (.A1(_09063_),
    .A2(_09064_),
    .B1(_09060_),
    .X(_09356_));
 sky130_fd_sc_hd__a21oi_4 _31700_ (.A1(_09353_),
    .A2(_09355_),
    .B1(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__clkbuf_4 _31701_ (.A(\pcpi_mul.rs1[26] ),
    .X(_09358_));
 sky130_fd_sc_hd__buf_4 _31702_ (.A(_09358_),
    .X(_09359_));
 sky130_fd_sc_hd__nand2_1 _31703_ (.A(_06636_),
    .B(_09075_),
    .Y(_09360_));
 sky130_fd_sc_hd__a21o_1 _31704_ (.A1(_05235_),
    .A2(_09359_),
    .B1(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__buf_4 _31705_ (.A(_09079_),
    .X(_09362_));
 sky130_fd_sc_hd__nand2_1 _31706_ (.A(_05163_),
    .B(_19848_),
    .Y(_09363_));
 sky130_fd_sc_hd__a21o_1 _31707_ (.A1(_06281_),
    .A2(_09362_),
    .B1(_09363_),
    .X(_09364_));
 sky130_fd_sc_hd__buf_6 _31708_ (.A(_08773_),
    .X(_09365_));
 sky130_fd_sc_hd__nand2_4 _31709_ (.A(_05807_),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__a21oi_4 _31710_ (.A1(_09361_),
    .A2(_09364_),
    .B1(_09366_),
    .Y(_09367_));
 sky130_fd_sc_hd__nand3_2 _31711_ (.A(_09361_),
    .B(_09364_),
    .C(_09366_),
    .Y(_09368_));
 sky130_vsdinv _31712_ (.A(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__nor2_4 _31713_ (.A(_09367_),
    .B(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__nand3_4 _31714_ (.A(_09353_),
    .B(_09356_),
    .C(_09355_),
    .Y(_09371_));
 sky130_fd_sc_hd__nand2_1 _31715_ (.A(_09370_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__nand3_2 _31716_ (.A(_09348_),
    .B(_09350_),
    .C(_09351_),
    .Y(_09373_));
 sky130_fd_sc_hd__a21oi_2 _31717_ (.A1(_09063_),
    .A2(_09064_),
    .B1(_09060_),
    .Y(_09374_));
 sky130_fd_sc_hd__o21ai_2 _31718_ (.A1(_09349_),
    .A2(_09354_),
    .B1(_09352_),
    .Y(_09375_));
 sky130_fd_sc_hd__nand3_4 _31719_ (.A(_09373_),
    .B(_09374_),
    .C(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__nand2_1 _31720_ (.A(_09371_),
    .B(_09376_),
    .Y(_09377_));
 sky130_fd_sc_hd__a21o_1 _31721_ (.A1(_09361_),
    .A2(_09364_),
    .B1(_09366_),
    .X(_09378_));
 sky130_fd_sc_hd__nand2_2 _31722_ (.A(_09378_),
    .B(_09368_),
    .Y(_09379_));
 sky130_fd_sc_hd__nand2_1 _31723_ (.A(_09377_),
    .B(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__nand2_1 _31724_ (.A(_09086_),
    .B(_09074_),
    .Y(_09381_));
 sky130_fd_sc_hd__nand2_1 _31725_ (.A(_09381_),
    .B(_09070_),
    .Y(_09382_));
 sky130_fd_sc_hd__o211ai_4 _31726_ (.A1(_09357_),
    .A2(_09372_),
    .B1(_09380_),
    .C1(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__a21boi_4 _31727_ (.A1(_09086_),
    .A2(_09074_),
    .B1_N(_09070_),
    .Y(_09384_));
 sky130_fd_sc_hd__nand2_2 _31728_ (.A(_09377_),
    .B(_09370_),
    .Y(_09385_));
 sky130_fd_sc_hd__nand3_4 _31729_ (.A(_09379_),
    .B(_09371_),
    .C(_09376_),
    .Y(_09386_));
 sky130_fd_sc_hd__o21ba_2 _31730_ (.A1(_09077_),
    .A2(_09080_),
    .B1_N(_09084_),
    .X(_09387_));
 sky130_fd_sc_hd__a31oi_4 _31731_ (.A1(_09384_),
    .A2(_09385_),
    .A3(_09386_),
    .B1(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__nand3_2 _31732_ (.A(_09384_),
    .B(_09385_),
    .C(_09386_),
    .Y(_09389_));
 sky130_fd_sc_hd__a21boi_4 _31733_ (.A1(_09383_),
    .A2(_09389_),
    .B1_N(_09387_),
    .Y(_09390_));
 sky130_fd_sc_hd__a21oi_4 _31734_ (.A1(_09383_),
    .A2(_09388_),
    .B1(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__nand2_1 _31735_ (.A(_09345_),
    .B(_09391_),
    .Y(_09392_));
 sky130_fd_sc_hd__and2_1 _31736_ (.A(_09388_),
    .B(_09383_),
    .X(_09393_));
 sky130_fd_sc_hd__o211ai_4 _31737_ (.A1(_09390_),
    .A2(_09393_),
    .B1(_09338_),
    .C1(_09344_),
    .Y(_09394_));
 sky130_fd_sc_hd__a21boi_2 _31738_ (.A1(_09185_),
    .A2(_09189_),
    .B1_N(_09182_),
    .Y(_09395_));
 sky130_fd_sc_hd__nand3_4 _31739_ (.A(_09392_),
    .B(_09394_),
    .C(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__nand2_1 _31740_ (.A(_09267_),
    .B(_09182_),
    .Y(_09397_));
 sky130_fd_sc_hd__o2bb2ai_2 _31741_ (.A1_N(_09338_),
    .A2_N(_09344_),
    .B1(_09393_),
    .B2(_09390_),
    .Y(_09398_));
 sky130_fd_sc_hd__nand3_2 _31742_ (.A(_09391_),
    .B(_09338_),
    .C(_09344_),
    .Y(_09399_));
 sky130_fd_sc_hd__nand3_4 _31743_ (.A(_09397_),
    .B(_09398_),
    .C(_09399_),
    .Y(_09400_));
 sky130_vsdinv _31744_ (.A(_09052_),
    .Y(_09401_));
 sky130_fd_sc_hd__a21o_2 _31745_ (.A1(_09103_),
    .A2(_09057_),
    .B1(_09401_),
    .X(_09402_));
 sky130_fd_sc_hd__a21oi_4 _31746_ (.A1(_09396_),
    .A2(_09400_),
    .B1(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__and2_1 _31747_ (.A(_09103_),
    .B(_09057_),
    .X(_09404_));
 sky130_fd_sc_hd__o211a_2 _31748_ (.A1(_09401_),
    .A2(_09404_),
    .B1(_09400_),
    .C1(_09396_),
    .X(_09405_));
 sky130_fd_sc_hd__nor2_4 _31749_ (.A(_09403_),
    .B(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__nand2_1 _31750_ (.A(_09245_),
    .B(_09242_),
    .Y(_09407_));
 sky130_fd_sc_hd__nand2_1 _31751_ (.A(_09255_),
    .B(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_1 _31752_ (.A(_09135_),
    .B(_09138_),
    .Y(_09409_));
 sky130_fd_sc_hd__a22oi_4 _31753_ (.A1(_06923_),
    .A2(_05643_),
    .B1(_08192_),
    .B2(_05976_),
    .Y(_09410_));
 sky130_fd_sc_hd__and4_2 _31754_ (.A(_19630_),
    .B(_19634_),
    .C(_06117_),
    .D(_19900_),
    .X(_09411_));
 sky130_fd_sc_hd__nand2_2 _31755_ (.A(\pcpi_mul.rs2[15] ),
    .B(_06287_),
    .Y(_09412_));
 sky130_fd_sc_hd__o21ai_2 _31756_ (.A1(_09410_),
    .A2(_09411_),
    .B1(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__nand2_1 _31757_ (.A(_19630_),
    .B(_05642_),
    .Y(_09414_));
 sky130_fd_sc_hd__nand3b_4 _31758_ (.A_N(_09414_),
    .B(_06988_),
    .C(_06648_),
    .Y(_09415_));
 sky130_vsdinv _31759_ (.A(_09412_),
    .Y(_09416_));
 sky130_fd_sc_hd__a22o_2 _31760_ (.A1(_07743_),
    .A2(_19900_),
    .B1(_06920_),
    .B2(_19897_),
    .X(_09417_));
 sky130_fd_sc_hd__nand3_2 _31761_ (.A(_09415_),
    .B(_09416_),
    .C(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__o21ai_2 _31762_ (.A1(_09212_),
    .A2(_09208_),
    .B1(_09214_),
    .Y(_09419_));
 sky130_fd_sc_hd__nand3_4 _31763_ (.A(_09413_),
    .B(_09418_),
    .C(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__o21ai_2 _31764_ (.A1(_09410_),
    .A2(_09411_),
    .B1(_09416_),
    .Y(_09421_));
 sky130_fd_sc_hd__nand3_4 _31765_ (.A(_09415_),
    .B(_09412_),
    .C(_09417_),
    .Y(_09422_));
 sky130_fd_sc_hd__a21oi_4 _31766_ (.A1(_09215_),
    .A2(_09216_),
    .B1(_09211_),
    .Y(_09423_));
 sky130_fd_sc_hd__nand3_4 _31767_ (.A(_09421_),
    .B(_09422_),
    .C(_09423_),
    .Y(_09424_));
 sky130_fd_sc_hd__nor2_2 _31768_ (.A(_09125_),
    .B(_09123_),
    .Y(_09425_));
 sky130_fd_sc_hd__o2bb2ai_4 _31769_ (.A1_N(_09420_),
    .A2_N(_09424_),
    .B1(_09121_),
    .B2(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__a21oi_2 _31770_ (.A1(_09129_),
    .A2(_09125_),
    .B1(_09123_),
    .Y(_09427_));
 sky130_fd_sc_hd__nand3b_4 _31771_ (.A_N(_09427_),
    .B(_09420_),
    .C(_09424_),
    .Y(_09428_));
 sky130_fd_sc_hd__a22oi_4 _31772_ (.A1(_09131_),
    .A2(_09409_),
    .B1(_09426_),
    .B2(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__a31oi_4 _31773_ (.A1(_09126_),
    .A2(_09128_),
    .A3(_09130_),
    .B1(_09138_),
    .Y(_09430_));
 sky130_vsdinv _31774_ (.A(_09135_),
    .Y(_09431_));
 sky130_fd_sc_hd__o211a_2 _31775_ (.A1(_09430_),
    .A2(_09431_),
    .B1(_09428_),
    .C1(_09426_),
    .X(_09432_));
 sky130_fd_sc_hd__a22oi_4 _31776_ (.A1(_06896_),
    .A2(_19891_),
    .B1(_06907_),
    .B2(_07064_),
    .Y(_09433_));
 sky130_fd_sc_hd__and4_1 _31777_ (.A(_06605_),
    .B(_19646_),
    .C(_06808_),
    .D(_19890_),
    .X(_09434_));
 sky130_fd_sc_hd__nand2_2 _31778_ (.A(_07223_),
    .B(_19883_),
    .Y(_09435_));
 sky130_vsdinv _31779_ (.A(_09435_),
    .Y(_09436_));
 sky130_fd_sc_hd__o21ai_2 _31780_ (.A1(_09433_),
    .A2(_09434_),
    .B1(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__nand2_1 _31781_ (.A(_06608_),
    .B(_06465_),
    .Y(_09438_));
 sky130_fd_sc_hd__buf_4 _31782_ (.A(_06168_),
    .X(_09439_));
 sky130_fd_sc_hd__nand3b_4 _31783_ (.A_N(_09438_),
    .B(_09439_),
    .C(_07327_),
    .Y(_09440_));
 sky130_fd_sc_hd__a22o_1 _31784_ (.A1(_06605_),
    .A2(_19890_),
    .B1(_06897_),
    .B2(_19887_),
    .X(_09441_));
 sky130_fd_sc_hd__nand3_4 _31785_ (.A(_09440_),
    .B(_09435_),
    .C(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__a21oi_4 _31786_ (.A1(_09151_),
    .A2(_09154_),
    .B1(_09149_),
    .Y(_09443_));
 sky130_fd_sc_hd__a21o_2 _31787_ (.A1(_09437_),
    .A2(_09442_),
    .B1(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__nand3_4 _31788_ (.A(_09437_),
    .B(_09442_),
    .C(_09443_),
    .Y(_09445_));
 sky130_fd_sc_hd__nand2_1 _31789_ (.A(_09444_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__a22oi_4 _31790_ (.A1(_06883_),
    .A2(_06799_),
    .B1(_06159_),
    .B2(_07056_),
    .Y(_09447_));
 sky130_fd_sc_hd__and4_1 _31791_ (.A(_06022_),
    .B(_06024_),
    .C(_06783_),
    .D(_06803_),
    .X(_09448_));
 sky130_fd_sc_hd__nand2_1 _31792_ (.A(_05731_),
    .B(_07067_),
    .Y(_09449_));
 sky130_vsdinv _31793_ (.A(_09449_),
    .Y(_09450_));
 sky130_fd_sc_hd__o21ai_1 _31794_ (.A1(_09447_),
    .A2(_09448_),
    .B1(_09450_),
    .Y(_09451_));
 sky130_fd_sc_hd__nand2_1 _31795_ (.A(_06326_),
    .B(_06654_),
    .Y(_09452_));
 sky130_fd_sc_hd__nand3b_4 _31796_ (.A_N(_09452_),
    .B(_19655_),
    .C(_19878_),
    .Y(_09453_));
 sky130_fd_sc_hd__a22o_1 _31797_ (.A1(_07893_),
    .A2(_08280_),
    .B1(_06335_),
    .B2(_07056_),
    .X(_09454_));
 sky130_fd_sc_hd__nand3_1 _31798_ (.A(_09453_),
    .B(_09449_),
    .C(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__nand2_2 _31799_ (.A(_09451_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__nand2_1 _31800_ (.A(_09446_),
    .B(_09456_),
    .Y(_09457_));
 sky130_vsdinv _31801_ (.A(_09456_),
    .Y(_09458_));
 sky130_fd_sc_hd__nand3_2 _31802_ (.A(_09458_),
    .B(_09444_),
    .C(_09445_),
    .Y(_09459_));
 sky130_fd_sc_hd__nand2_4 _31803_ (.A(_09457_),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__o21ai_4 _31804_ (.A1(_09429_),
    .A2(_09432_),
    .B1(_09460_),
    .Y(_09461_));
 sky130_fd_sc_hd__nand2_2 _31805_ (.A(_09140_),
    .B(_09135_),
    .Y(_09462_));
 sky130_fd_sc_hd__a21o_2 _31806_ (.A1(_09426_),
    .A2(_09428_),
    .B1(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__nand2_1 _31807_ (.A(_09446_),
    .B(_09458_),
    .Y(_09464_));
 sky130_fd_sc_hd__nand3_1 _31808_ (.A(_09444_),
    .B(_09456_),
    .C(_09445_),
    .Y(_09465_));
 sky130_fd_sc_hd__nand2_2 _31809_ (.A(_09464_),
    .B(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand3_4 _31810_ (.A(_09462_),
    .B(_09428_),
    .C(_09426_),
    .Y(_09467_));
 sky130_fd_sc_hd__nand3_4 _31811_ (.A(_09463_),
    .B(_09466_),
    .C(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__nand3_4 _31812_ (.A(_09461_),
    .B(_09241_),
    .C(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__o21ai_2 _31813_ (.A1(_09429_),
    .A2(_09432_),
    .B1(_09466_),
    .Y(_09470_));
 sky130_fd_sc_hd__nand3_4 _31814_ (.A(_09463_),
    .B(_09460_),
    .C(_09467_),
    .Y(_09471_));
 sky130_fd_sc_hd__nand3_4 _31815_ (.A(_09470_),
    .B(_09249_),
    .C(_09471_),
    .Y(_09472_));
 sky130_fd_sc_hd__nor2_4 _31816_ (.A(_09179_),
    .B(_09144_),
    .Y(_09473_));
 sky130_fd_sc_hd__nor2_4 _31817_ (.A(_09141_),
    .B(_09473_),
    .Y(_09474_));
 sky130_fd_sc_hd__a21oi_4 _31818_ (.A1(_09469_),
    .A2(_09472_),
    .B1(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__nor2_2 _31819_ (.A(_09174_),
    .B(_09141_),
    .Y(_09476_));
 sky130_fd_sc_hd__o211a_1 _31820_ (.A1(_09144_),
    .A2(_09476_),
    .B1(_09469_),
    .C1(_09472_),
    .X(_09477_));
 sky130_fd_sc_hd__nand2_4 _31821_ (.A(_19595_),
    .B(_05105_),
    .Y(_09478_));
 sky130_fd_sc_hd__nand2_4 _31822_ (.A(_08945_),
    .B(_05229_),
    .Y(_09479_));
 sky130_fd_sc_hd__or2_2 _31823_ (.A(_09478_),
    .B(_09479_),
    .X(_09480_));
 sky130_fd_sc_hd__nand2_2 _31824_ (.A(\pcpi_mul.rs2[24] ),
    .B(_05263_),
    .Y(_09481_));
 sky130_fd_sc_hd__nand2_4 _31825_ (.A(_09478_),
    .B(_09479_),
    .Y(_09482_));
 sky130_fd_sc_hd__nand3_4 _31826_ (.A(_09480_),
    .B(_09481_),
    .C(_09482_),
    .Y(_09483_));
 sky130_fd_sc_hd__a21oi_4 _31827_ (.A1(_09233_),
    .A2(_09235_),
    .B1(_09231_),
    .Y(_09484_));
 sky130_fd_sc_hd__buf_8 _31828_ (.A(_09229_),
    .X(_09485_));
 sky130_fd_sc_hd__a22oi_4 _31829_ (.A1(_09485_),
    .A2(_07759_),
    .B1(_19600_),
    .B2(_05121_),
    .Y(_09486_));
 sky130_fd_sc_hd__nor2_8 _31830_ (.A(_09478_),
    .B(_09479_),
    .Y(_09487_));
 sky130_vsdinv _31831_ (.A(_09481_),
    .Y(_09488_));
 sky130_fd_sc_hd__o21ai_4 _31832_ (.A1(_09486_),
    .A2(_09487_),
    .B1(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__nand2_2 _31833_ (.A(_19592_),
    .B(_19934_),
    .Y(_09490_));
 sky130_fd_sc_hd__a31oi_4 _31834_ (.A1(_09483_),
    .A2(_09484_),
    .A3(_09489_),
    .B1(_09490_),
    .Y(_09491_));
 sky130_fd_sc_hd__o21ai_2 _31835_ (.A1(_09486_),
    .A2(_09487_),
    .B1(_09481_),
    .Y(_09492_));
 sky130_fd_sc_hd__nand3_2 _31836_ (.A(_09480_),
    .B(_09488_),
    .C(_09482_),
    .Y(_09493_));
 sky130_fd_sc_hd__nand3b_4 _31837_ (.A_N(_09484_),
    .B(_09492_),
    .C(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__nand2_1 _31838_ (.A(_09491_),
    .B(_09494_),
    .Y(_09495_));
 sky130_vsdinv _31839_ (.A(_09495_),
    .Y(_09496_));
 sky130_fd_sc_hd__nand3_2 _31840_ (.A(_09483_),
    .B(_09484_),
    .C(_09489_),
    .Y(_09497_));
 sky130_fd_sc_hd__a21boi_4 _31841_ (.A1(_09494_),
    .A2(_09497_),
    .B1_N(_09490_),
    .Y(_09498_));
 sky130_fd_sc_hd__nand3_4 _31842_ (.A(_19620_),
    .B(_19624_),
    .C(_05480_),
    .Y(_09499_));
 sky130_fd_sc_hd__nor2_8 _31843_ (.A(_05663_),
    .B(_09499_),
    .Y(_09500_));
 sky130_fd_sc_hd__a22o_1 _31844_ (.A1(_07933_),
    .A2(_05488_),
    .B1(_07824_),
    .B2(_19906_),
    .X(_09501_));
 sky130_fd_sc_hd__nand2_4 _31845_ (.A(\pcpi_mul.rs2[18] ),
    .B(_19903_),
    .Y(_09502_));
 sky130_fd_sc_hd__nand3b_2 _31846_ (.A_N(_09500_),
    .B(_09501_),
    .C(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__a22oi_4 _31847_ (.A1(_07933_),
    .A2(_05769_),
    .B1(_07824_),
    .B2(_05464_),
    .Y(_09504_));
 sky130_vsdinv _31848_ (.A(_09502_),
    .Y(_09505_));
 sky130_fd_sc_hd__o21ai_2 _31849_ (.A1(_09504_),
    .A2(_09500_),
    .B1(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__nand2_4 _31850_ (.A(_09503_),
    .B(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__a22oi_4 _31851_ (.A1(_09191_),
    .A2(_05173_),
    .B1(_08154_),
    .B2(_05377_),
    .Y(_09508_));
 sky130_fd_sc_hd__clkinv_8 _31852_ (.A(\pcpi_mul.rs1[5] ),
    .Y(_09509_));
 sky130_fd_sc_hd__nand3_4 _31853_ (.A(_19606_),
    .B(_19610_),
    .C(_05172_),
    .Y(_09510_));
 sky130_fd_sc_hd__nor2_4 _31854_ (.A(_09509_),
    .B(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__nand2_4 _31855_ (.A(\pcpi_mul.rs2[21] ),
    .B(_19912_),
    .Y(_09512_));
 sky130_vsdinv _31856_ (.A(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__o21ai_2 _31857_ (.A1(_09508_),
    .A2(_09511_),
    .B1(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__a21oi_2 _31858_ (.A1(_09199_),
    .A2(_09200_),
    .B1(_09195_),
    .Y(_09515_));
 sky130_fd_sc_hd__clkbuf_4 _31859_ (.A(\pcpi_mul.rs2[22] ),
    .X(_09516_));
 sky130_fd_sc_hd__a22o_2 _31860_ (.A1(_09191_),
    .A2(_05173_),
    .B1(_09516_),
    .B2(_19916_),
    .X(_09517_));
 sky130_fd_sc_hd__o211ai_4 _31861_ (.A1(_09509_),
    .A2(_09510_),
    .B1(_09512_),
    .C1(_09517_),
    .Y(_09518_));
 sky130_fd_sc_hd__nand3_4 _31862_ (.A(_09514_),
    .B(_09515_),
    .C(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__o21ai_2 _31863_ (.A1(_09508_),
    .A2(_09511_),
    .B1(_09512_),
    .Y(_09520_));
 sky130_fd_sc_hd__o21ai_2 _31864_ (.A1(_09196_),
    .A2(_09192_),
    .B1(_09198_),
    .Y(_09521_));
 sky130_fd_sc_hd__o211ai_4 _31865_ (.A1(_09509_),
    .A2(_09510_),
    .B1(_09513_),
    .C1(_09517_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand3_4 _31866_ (.A(_09520_),
    .B(_09521_),
    .C(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__nand3_4 _31867_ (.A(_09507_),
    .B(_09519_),
    .C(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__o21a_1 _31868_ (.A1(_09504_),
    .A2(_09500_),
    .B1(_09502_),
    .X(_09525_));
 sky130_fd_sc_hd__nor3_4 _31869_ (.A(_09502_),
    .B(_09504_),
    .C(_09500_),
    .Y(_09526_));
 sky130_fd_sc_hd__o2bb2ai_4 _31870_ (.A1_N(_09523_),
    .A2_N(_09519_),
    .B1(_09525_),
    .B2(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__o2bb2ai_4 _31871_ (.A1_N(_09524_),
    .A2_N(_09527_),
    .B1(_09226_),
    .B2(_09237_),
    .Y(_09528_));
 sky130_fd_sc_hd__nand3_4 _31872_ (.A(_09527_),
    .B(_09238_),
    .C(_09524_),
    .Y(_09529_));
 sky130_fd_sc_hd__nand2_4 _31873_ (.A(_09247_),
    .B(_09203_),
    .Y(_09530_));
 sky130_fd_sc_hd__a21oi_4 _31874_ (.A1(_09528_),
    .A2(_09529_),
    .B1(_09530_),
    .Y(_09531_));
 sky130_vsdinv _31875_ (.A(_09530_),
    .Y(_09532_));
 sky130_fd_sc_hd__a21oi_4 _31876_ (.A1(_09527_),
    .A2(_09524_),
    .B1(_09238_),
    .Y(_09533_));
 sky130_fd_sc_hd__nand2_1 _31877_ (.A(_09507_),
    .B(_09523_),
    .Y(_09534_));
 sky130_vsdinv _31878_ (.A(_09519_),
    .Y(_09535_));
 sky130_fd_sc_hd__o211a_4 _31879_ (.A1(_09534_),
    .A2(_09535_),
    .B1(_09238_),
    .C1(_09527_),
    .X(_09536_));
 sky130_fd_sc_hd__nor3_4 _31880_ (.A(_09532_),
    .B(_09533_),
    .C(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__o22ai_4 _31881_ (.A1(_09496_),
    .A2(_09498_),
    .B1(_09531_),
    .B2(_09537_),
    .Y(_09538_));
 sky130_fd_sc_hd__o21ai_2 _31882_ (.A1(_09533_),
    .A2(_09536_),
    .B1(_09532_),
    .Y(_09539_));
 sky130_fd_sc_hd__nand3_4 _31883_ (.A(_09528_),
    .B(_09529_),
    .C(_09530_),
    .Y(_09540_));
 sky130_fd_sc_hd__nor2_2 _31884_ (.A(_09498_),
    .B(_09496_),
    .Y(_09541_));
 sky130_fd_sc_hd__nand3_4 _31885_ (.A(_09539_),
    .B(_09540_),
    .C(_09541_),
    .Y(_09542_));
 sky130_vsdinv _31886_ (.A(_09242_),
    .Y(_09543_));
 sky130_fd_sc_hd__a21oi_4 _31887_ (.A1(_09538_),
    .A2(_09542_),
    .B1(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__nand2_1 _31888_ (.A(_09539_),
    .B(_09541_),
    .Y(_09545_));
 sky130_fd_sc_hd__o211a_2 _31889_ (.A1(_09537_),
    .A2(_09545_),
    .B1(_09543_),
    .C1(_09538_),
    .X(_09546_));
 sky130_fd_sc_hd__o22ai_4 _31890_ (.A1(_09475_),
    .A2(_09477_),
    .B1(_09544_),
    .B2(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__and3_2 _31891_ (.A(_09470_),
    .B(_09471_),
    .C(_09249_),
    .X(_09548_));
 sky130_fd_sc_hd__nand2_4 _31892_ (.A(_09469_),
    .B(_09474_),
    .Y(_09549_));
 sky130_fd_sc_hd__o2bb2ai_4 _31893_ (.A1_N(_09469_),
    .A2_N(_09472_),
    .B1(_09141_),
    .B2(_09473_),
    .Y(_09550_));
 sky130_fd_sc_hd__nand3_4 _31894_ (.A(_09538_),
    .B(_09543_),
    .C(_09542_),
    .Y(_09551_));
 sky130_fd_sc_hd__nand2_1 _31895_ (.A(_09538_),
    .B(_09542_),
    .Y(_09552_));
 sky130_fd_sc_hd__nand2_4 _31896_ (.A(_09552_),
    .B(_09242_),
    .Y(_09553_));
 sky130_fd_sc_hd__o2111ai_4 _31897_ (.A1(_09548_),
    .A2(_09549_),
    .B1(_09550_),
    .C1(_09551_),
    .D1(_09553_),
    .Y(_09554_));
 sky130_fd_sc_hd__nand3_4 _31898_ (.A(_09408_),
    .B(_09547_),
    .C(_09554_),
    .Y(_09555_));
 sky130_fd_sc_hd__nor2_2 _31899_ (.A(_09144_),
    .B(_09476_),
    .Y(_09556_));
 sky130_fd_sc_hd__a31oi_4 _31900_ (.A1(_09241_),
    .A2(_09461_),
    .A3(_09468_),
    .B1(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__a21oi_4 _31901_ (.A1(_09472_),
    .A2(_09557_),
    .B1(_09475_),
    .Y(_09558_));
 sky130_fd_sc_hd__o21ai_2 _31902_ (.A1(_09544_),
    .A2(_09546_),
    .B1(_09558_),
    .Y(_09559_));
 sky130_vsdinv _31903_ (.A(_09407_),
    .Y(_09560_));
 sky130_fd_sc_hd__a31oi_4 _31904_ (.A1(_09253_),
    .A2(_09188_),
    .A3(_09190_),
    .B1(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__o21ai_4 _31905_ (.A1(_09548_),
    .A2(_09549_),
    .B1(_09550_),
    .Y(_09562_));
 sky130_fd_sc_hd__nand3_4 _31906_ (.A(_09562_),
    .B(_09553_),
    .C(_09551_),
    .Y(_09563_));
 sky130_fd_sc_hd__nand3_4 _31907_ (.A(_09559_),
    .B(_09561_),
    .C(_09563_),
    .Y(_09564_));
 sky130_fd_sc_hd__nand3_2 _31908_ (.A(_09406_),
    .B(_09555_),
    .C(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand2_2 _31909_ (.A(_09564_),
    .B(_09555_),
    .Y(_09566_));
 sky130_fd_sc_hd__o21ai_2 _31910_ (.A1(_09403_),
    .A2(_09405_),
    .B1(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand3_4 _31911_ (.A(_09306_),
    .B(_09565_),
    .C(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__a31oi_4 _31912_ (.A1(_09119_),
    .A2(_09270_),
    .A3(_09116_),
    .B1(_09261_),
    .Y(_09569_));
 sky130_fd_sc_hd__nand2_4 _31913_ (.A(_09406_),
    .B(_09566_),
    .Y(_09570_));
 sky130_fd_sc_hd__o211ai_4 _31914_ (.A1(_09403_),
    .A2(_09405_),
    .B1(_09555_),
    .C1(_09564_),
    .Y(_09571_));
 sky130_fd_sc_hd__nand3_4 _31915_ (.A(_09569_),
    .B(_09570_),
    .C(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__nand2_2 _31916_ (.A(_09568_),
    .B(_09572_),
    .Y(_09573_));
 sky130_fd_sc_hd__and2_1 _31917_ (.A(_09097_),
    .B(_09092_),
    .X(_09574_));
 sky130_fd_sc_hd__a21o_4 _31918_ (.A1(_09264_),
    .A2(_09113_),
    .B1(_09574_),
    .X(_09575_));
 sky130_fd_sc_hd__nand3_4 _31919_ (.A(_09264_),
    .B(_09113_),
    .C(_09574_),
    .Y(_09576_));
 sky130_fd_sc_hd__nand2_4 _31920_ (.A(_09575_),
    .B(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__nand2_1 _31921_ (.A(_09573_),
    .B(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__o21ai_2 _31922_ (.A1(_09288_),
    .A2(_09275_),
    .B1(_09282_),
    .Y(_09579_));
 sky130_fd_sc_hd__a31oi_4 _31923_ (.A1(_09569_),
    .A2(_09570_),
    .A3(_09571_),
    .B1(_09577_),
    .Y(_09580_));
 sky130_fd_sc_hd__nand2_1 _31924_ (.A(_09580_),
    .B(_09568_),
    .Y(_09581_));
 sky130_fd_sc_hd__nand3_4 _31925_ (.A(_09578_),
    .B(_09579_),
    .C(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__a21oi_4 _31926_ (.A1(_09281_),
    .A2(_09283_),
    .B1(_09278_),
    .Y(_09583_));
 sky130_fd_sc_hd__nand3_4 _31927_ (.A(_09568_),
    .B(_09572_),
    .C(_09577_),
    .Y(_09584_));
 sky130_fd_sc_hd__and2_1 _31928_ (.A(_09575_),
    .B(_09576_),
    .X(_09585_));
 sky130_fd_sc_hd__nand2_4 _31929_ (.A(_09573_),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__nand3_4 _31930_ (.A(_09583_),
    .B(_09584_),
    .C(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__and2_1 _31931_ (.A(_08975_),
    .B(_08832_),
    .X(_09588_));
 sky130_fd_sc_hd__o2bb2ai_2 _31932_ (.A1_N(_09582_),
    .A2_N(_09587_),
    .B1(_09588_),
    .B2(_09015_),
    .Y(_09589_));
 sky130_fd_sc_hd__nand3_4 _31933_ (.A(_09587_),
    .B(_09582_),
    .C(_09016_),
    .Y(_09590_));
 sky130_fd_sc_hd__nand2_1 _31934_ (.A(_09298_),
    .B(_09285_),
    .Y(_09591_));
 sky130_fd_sc_hd__a21oi_4 _31935_ (.A1(_09589_),
    .A2(_09590_),
    .B1(_09591_),
    .Y(_09592_));
 sky130_vsdinv _31936_ (.A(_08986_),
    .Y(_09593_));
 sky130_fd_sc_hd__a31oi_1 _31937_ (.A1(_09286_),
    .A2(_09289_),
    .A3(_09287_),
    .B1(_09593_),
    .Y(_09594_));
 sky130_fd_sc_hd__o211a_2 _31938_ (.A1(_09297_),
    .A2(_09594_),
    .B1(_09590_),
    .C1(_09589_),
    .X(_09595_));
 sky130_fd_sc_hd__nor2_8 _31939_ (.A(_09592_),
    .B(_09595_),
    .Y(_09596_));
 sky130_vsdinv _31940_ (.A(_09299_),
    .Y(_09597_));
 sky130_fd_sc_hd__o21ai_4 _31941_ (.A1(_09296_),
    .A2(_09304_),
    .B1(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__xor2_4 _31942_ (.A(_09596_),
    .B(_09598_),
    .X(_02646_));
 sky130_fd_sc_hd__nor2_2 _31943_ (.A(_09432_),
    .B(_09460_),
    .Y(_09599_));
 sky130_fd_sc_hd__nand2_2 _31944_ (.A(_09532_),
    .B(_09529_),
    .Y(_09600_));
 sky130_fd_sc_hd__a22oi_4 _31945_ (.A1(_06022_),
    .A2(_06783_),
    .B1(_05736_),
    .B2(_07067_),
    .Y(_09601_));
 sky130_fd_sc_hd__and4_1 _31946_ (.A(_06401_),
    .B(_06158_),
    .C(_07554_),
    .D(_07050_),
    .X(_09602_));
 sky130_fd_sc_hd__nand2_1 _31947_ (.A(_19658_),
    .B(_08061_),
    .Y(_09603_));
 sky130_vsdinv _31948_ (.A(_09603_),
    .Y(_09604_));
 sky130_fd_sc_hd__o21ai_1 _31949_ (.A1(_09601_),
    .A2(_09602_),
    .B1(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__nand2_1 _31950_ (.A(_19651_),
    .B(_07050_),
    .Y(_09606_));
 sky130_fd_sc_hd__buf_6 _31951_ (.A(_07554_),
    .X(_09607_));
 sky130_fd_sc_hd__nand3b_2 _31952_ (.A_N(_09606_),
    .B(_06884_),
    .C(_09607_),
    .Y(_09608_));
 sky130_fd_sc_hd__a22o_1 _31953_ (.A1(_06326_),
    .A2(_19877_),
    .B1(_19654_),
    .B2(_19873_),
    .X(_09609_));
 sky130_fd_sc_hd__nand3_1 _31954_ (.A(_09608_),
    .B(_09609_),
    .C(_09603_),
    .Y(_09610_));
 sky130_fd_sc_hd__nand2_1 _31955_ (.A(_09605_),
    .B(_09610_),
    .Y(_09611_));
 sky130_vsdinv _31956_ (.A(_09611_),
    .Y(_09612_));
 sky130_fd_sc_hd__a21oi_2 _31957_ (.A1(_09441_),
    .A2(_09436_),
    .B1(_09434_),
    .Y(_09613_));
 sky130_fd_sc_hd__a22oi_4 _31958_ (.A1(_06608_),
    .A2(_07642_),
    .B1(_06610_),
    .B2(_06634_),
    .Y(_09614_));
 sky130_fd_sc_hd__and4_4 _31959_ (.A(_19643_),
    .B(_06167_),
    .C(\pcpi_mul.rs1[15] ),
    .D(_19886_),
    .X(_09615_));
 sky130_fd_sc_hd__nand2_2 _31960_ (.A(_07223_),
    .B(_06798_),
    .Y(_09616_));
 sky130_fd_sc_hd__o21ai_2 _31961_ (.A1(_09614_),
    .A2(_09615_),
    .B1(_09616_),
    .Y(_09617_));
 sky130_vsdinv _31962_ (.A(_09616_),
    .Y(_09618_));
 sky130_fd_sc_hd__a22o_2 _31963_ (.A1(_08219_),
    .A2(_06464_),
    .B1(_06168_),
    .B2(_06443_),
    .X(_09619_));
 sky130_fd_sc_hd__nand3b_4 _31964_ (.A_N(_09615_),
    .B(_09618_),
    .C(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__nand3b_4 _31965_ (.A_N(_09613_),
    .B(_09617_),
    .C(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__nand3b_1 _31966_ (.A_N(_09615_),
    .B(_09616_),
    .C(_09619_),
    .Y(_09622_));
 sky130_fd_sc_hd__o21ai_1 _31967_ (.A1(_09614_),
    .A2(_09615_),
    .B1(_09618_),
    .Y(_09623_));
 sky130_fd_sc_hd__nand3_2 _31968_ (.A(_09622_),
    .B(_09613_),
    .C(_09623_),
    .Y(_09624_));
 sky130_fd_sc_hd__nand2_1 _31969_ (.A(_09621_),
    .B(_09624_),
    .Y(_09625_));
 sky130_fd_sc_hd__nor2_2 _31970_ (.A(_09612_),
    .B(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__and2_1 _31971_ (.A(_09625_),
    .B(_09612_),
    .X(_09627_));
 sky130_fd_sc_hd__nand2_1 _31972_ (.A(_09420_),
    .B(_09427_),
    .Y(_09628_));
 sky130_fd_sc_hd__a22oi_4 _31973_ (.A1(_06923_),
    .A2(_05976_),
    .B1(_08192_),
    .B2(_06115_),
    .Y(_09629_));
 sky130_fd_sc_hd__and4_1 _31974_ (.A(_07743_),
    .B(_19634_),
    .C(_06287_),
    .D(_19897_),
    .X(_09630_));
 sky130_fd_sc_hd__nand2_4 _31975_ (.A(_19640_),
    .B(_06282_),
    .Y(_09631_));
 sky130_vsdinv _31976_ (.A(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__o21ai_2 _31977_ (.A1(_09629_),
    .A2(_09630_),
    .B1(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__a21oi_4 _31978_ (.A1(_09501_),
    .A2(_09505_),
    .B1(_09500_),
    .Y(_09634_));
 sky130_fd_sc_hd__nand2_1 _31979_ (.A(_19630_),
    .B(_06117_),
    .Y(_09635_));
 sky130_fd_sc_hd__nand3b_4 _31980_ (.A_N(_09635_),
    .B(_07428_),
    .C(_07502_),
    .Y(_09636_));
 sky130_fd_sc_hd__a22o_1 _31981_ (.A1(_07923_),
    .A2(_05976_),
    .B1(_08192_),
    .B2(_06115_),
    .X(_09637_));
 sky130_fd_sc_hd__nand3_4 _31982_ (.A(_09636_),
    .B(_09631_),
    .C(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__nand3_4 _31983_ (.A(_09633_),
    .B(_09634_),
    .C(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__o21ai_2 _31984_ (.A1(_09629_),
    .A2(_09630_),
    .B1(_09631_),
    .Y(_09640_));
 sky130_fd_sc_hd__nand3_2 _31985_ (.A(_09636_),
    .B(_09632_),
    .C(_09637_),
    .Y(_09641_));
 sky130_fd_sc_hd__o22ai_4 _31986_ (.A1(net449),
    .A2(_09499_),
    .B1(_09502_),
    .B2(_09504_),
    .Y(_09642_));
 sky130_fd_sc_hd__nand3_4 _31987_ (.A(_09640_),
    .B(_09641_),
    .C(_09642_),
    .Y(_09643_));
 sky130_fd_sc_hd__nand2_1 _31988_ (.A(_09639_),
    .B(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__a21oi_4 _31989_ (.A1(_09417_),
    .A2(_09416_),
    .B1(_09411_),
    .Y(_09645_));
 sky130_fd_sc_hd__nand2_4 _31990_ (.A(_09644_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__nand3b_4 _31991_ (.A_N(_09645_),
    .B(_09639_),
    .C(_09643_),
    .Y(_09647_));
 sky130_fd_sc_hd__a22oi_4 _31992_ (.A1(_09424_),
    .A2(_09628_),
    .B1(_09646_),
    .B2(_09647_),
    .Y(_09648_));
 sky130_vsdinv _31993_ (.A(_09420_),
    .Y(_09649_));
 sky130_fd_sc_hd__a31oi_1 _31994_ (.A1(_09421_),
    .A2(_09422_),
    .A3(_09423_),
    .B1(_09427_),
    .Y(_09650_));
 sky130_fd_sc_hd__o211a_1 _31995_ (.A1(_09649_),
    .A2(_09650_),
    .B1(_09647_),
    .C1(_09646_),
    .X(_09651_));
 sky130_fd_sc_hd__o22ai_4 _31996_ (.A1(_09626_),
    .A2(_09627_),
    .B1(_09648_),
    .B2(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__nand2_2 _31997_ (.A(_09428_),
    .B(_09420_),
    .Y(_09653_));
 sky130_fd_sc_hd__a21o_1 _31998_ (.A1(_09646_),
    .A2(_09647_),
    .B1(_09653_),
    .X(_09654_));
 sky130_fd_sc_hd__nand3_4 _31999_ (.A(_09653_),
    .B(_09647_),
    .C(_09646_),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_1 _32000_ (.A(_09625_),
    .B(_09611_),
    .Y(_09656_));
 sky130_fd_sc_hd__nand3_1 _32001_ (.A(_09612_),
    .B(_09621_),
    .C(_09624_),
    .Y(_09657_));
 sky130_fd_sc_hd__nand2_1 _32002_ (.A(_09656_),
    .B(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__nand3_4 _32003_ (.A(_09654_),
    .B(_09655_),
    .C(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__a22oi_4 _32004_ (.A1(_09528_),
    .A2(_09600_),
    .B1(_09652_),
    .B2(_09659_),
    .Y(_09660_));
 sky130_fd_sc_hd__nor2_2 _32005_ (.A(_09532_),
    .B(_09533_),
    .Y(_09661_));
 sky130_fd_sc_hd__o211a_2 _32006_ (.A1(_09536_),
    .A2(_09661_),
    .B1(_09659_),
    .C1(_09652_),
    .X(_09662_));
 sky130_fd_sc_hd__o22ai_4 _32007_ (.A1(_09429_),
    .A2(_09599_),
    .B1(_09660_),
    .B2(_09662_),
    .Y(_09663_));
 sky130_fd_sc_hd__buf_2 _32008_ (.A(_09663_),
    .X(_09664_));
 sky130_vsdinv _32009_ (.A(_09600_),
    .Y(_09665_));
 sky130_fd_sc_hd__o2bb2ai_2 _32010_ (.A1_N(_09659_),
    .A2_N(_09652_),
    .B1(_09533_),
    .B2(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__o211ai_4 _32011_ (.A1(_09536_),
    .A2(_09661_),
    .B1(_09659_),
    .C1(_09652_),
    .Y(_09667_));
 sky130_fd_sc_hd__nand2_1 _32012_ (.A(_09463_),
    .B(_09460_),
    .Y(_09668_));
 sky130_fd_sc_hd__nand2_1 _32013_ (.A(_09668_),
    .B(_09467_),
    .Y(_09669_));
 sky130_fd_sc_hd__nand3_2 _32014_ (.A(_09666_),
    .B(_09667_),
    .C(_09669_),
    .Y(_09670_));
 sky130_fd_sc_hd__clkbuf_4 _32015_ (.A(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__nand2_1 _32016_ (.A(_09664_),
    .B(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__a22oi_4 _32017_ (.A1(_08152_),
    .A2(_05208_),
    .B1(_19611_),
    .B2(_05486_),
    .Y(_09673_));
 sky130_fd_sc_hd__nand3_4 _32018_ (.A(_08539_),
    .B(_09516_),
    .C(_05271_),
    .Y(_09674_));
 sky130_fd_sc_hd__nor2_2 _32019_ (.A(_05278_),
    .B(_09674_),
    .Y(_09675_));
 sky130_fd_sc_hd__nand2_4 _32020_ (.A(_08545_),
    .B(_05488_),
    .Y(_09676_));
 sky130_fd_sc_hd__o21ai_2 _32021_ (.A1(_09673_),
    .A2(_09675_),
    .B1(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__o22ai_4 _32022_ (.A1(_09509_),
    .A2(_09510_),
    .B1(_09512_),
    .B2(_09508_),
    .Y(_09678_));
 sky130_vsdinv _32023_ (.A(_09676_),
    .Y(_09679_));
 sky130_fd_sc_hd__buf_2 _32024_ (.A(_19610_),
    .X(_09680_));
 sky130_fd_sc_hd__a22o_2 _32025_ (.A1(_19607_),
    .A2(_05553_),
    .B1(_09680_),
    .B2(_05291_),
    .X(_09681_));
 sky130_fd_sc_hd__o211ai_4 _32026_ (.A1(net451),
    .A2(_09674_),
    .B1(_09679_),
    .C1(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__nand3_4 _32027_ (.A(_09677_),
    .B(_09678_),
    .C(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__o21ai_2 _32028_ (.A1(_09673_),
    .A2(_09675_),
    .B1(_09679_),
    .Y(_09684_));
 sky130_fd_sc_hd__a21oi_2 _32029_ (.A1(_09517_),
    .A2(_09513_),
    .B1(_09511_),
    .Y(_09685_));
 sky130_fd_sc_hd__o211ai_4 _32030_ (.A1(net451),
    .A2(_09674_),
    .B1(_09676_),
    .C1(_09681_),
    .Y(_09686_));
 sky130_fd_sc_hd__nand3_4 _32031_ (.A(_09684_),
    .B(_09685_),
    .C(_09686_),
    .Y(_09687_));
 sky130_fd_sc_hd__nand2_1 _32032_ (.A(_07822_),
    .B(_05464_),
    .Y(_09688_));
 sky130_fd_sc_hd__nand3b_4 _32033_ (.A_N(_09688_),
    .B(_08172_),
    .C(_06494_),
    .Y(_09689_));
 sky130_fd_sc_hd__a22o_2 _32034_ (.A1(_19621_),
    .A2(_05672_),
    .B1(_08174_),
    .B2(_06264_),
    .X(_09690_));
 sky130_fd_sc_hd__nand2_2 _32035_ (.A(_07481_),
    .B(_05643_),
    .Y(_09691_));
 sky130_vsdinv _32036_ (.A(_09691_),
    .Y(_09692_));
 sky130_fd_sc_hd__a21oi_2 _32037_ (.A1(_09689_),
    .A2(_09690_),
    .B1(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__and3_1 _32038_ (.A(_09689_),
    .B(_09692_),
    .C(_09690_),
    .X(_09694_));
 sky130_fd_sc_hd__o2bb2ai_4 _32039_ (.A1_N(_09683_),
    .A2_N(_09687_),
    .B1(_09693_),
    .B2(_09694_),
    .Y(_09695_));
 sky130_fd_sc_hd__a22oi_4 _32040_ (.A1(_07486_),
    .A2(_05672_),
    .B1(_08172_),
    .B2(_19904_),
    .Y(_09696_));
 sky130_fd_sc_hd__and4_1 _32041_ (.A(_19621_),
    .B(_07827_),
    .C(_05796_),
    .D(_05464_),
    .X(_09697_));
 sky130_fd_sc_hd__o21ai_1 _32042_ (.A1(_09696_),
    .A2(_09697_),
    .B1(_09692_),
    .Y(_09698_));
 sky130_fd_sc_hd__nand3_2 _32043_ (.A(_09689_),
    .B(_09691_),
    .C(_09690_),
    .Y(_09699_));
 sky130_fd_sc_hd__nand2_2 _32044_ (.A(_09698_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__nand3_4 _32045_ (.A(_09687_),
    .B(_09683_),
    .C(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__a21oi_4 _32046_ (.A1(_09483_),
    .A2(_09489_),
    .B1(_09484_),
    .Y(_09702_));
 sky130_fd_sc_hd__a21oi_4 _32047_ (.A1(_09695_),
    .A2(_09701_),
    .B1(_09702_),
    .Y(_09703_));
 sky130_fd_sc_hd__and3_2 _32048_ (.A(_09695_),
    .B(_09702_),
    .C(_09701_),
    .X(_09704_));
 sky130_fd_sc_hd__nand2_4 _32049_ (.A(_09524_),
    .B(_09523_),
    .Y(_09705_));
 sky130_vsdinv _32050_ (.A(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__o21ai_4 _32051_ (.A1(_09703_),
    .A2(_09704_),
    .B1(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__nand2_2 _32052_ (.A(_19586_),
    .B(_19932_),
    .Y(_09708_));
 sky130_fd_sc_hd__nand2_2 _32053_ (.A(\pcpi_mul.rs2[27] ),
    .B(_05122_),
    .Y(_09709_));
 sky130_fd_sc_hd__nor2_8 _32054_ (.A(_09708_),
    .B(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__and2_2 _32055_ (.A(_09708_),
    .B(_09709_),
    .X(_09711_));
 sky130_fd_sc_hd__nor2_8 _32056_ (.A(_09710_),
    .B(_09711_),
    .Y(_09712_));
 sky130_vsdinv _32057_ (.A(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__nand2_2 _32058_ (.A(_09229_),
    .B(_07828_),
    .Y(_09714_));
 sky130_fd_sc_hd__nand2_2 _32059_ (.A(_19599_),
    .B(_05695_),
    .Y(_09715_));
 sky130_fd_sc_hd__or2_2 _32060_ (.A(_09714_),
    .B(_09715_),
    .X(_09716_));
 sky130_fd_sc_hd__nand2_2 _32061_ (.A(_09714_),
    .B(_09715_),
    .Y(_09717_));
 sky130_fd_sc_hd__nand2_2 _32062_ (.A(_19602_),
    .B(_05272_),
    .Y(_09718_));
 sky130_vsdinv _32063_ (.A(_09718_),
    .Y(_09719_));
 sky130_fd_sc_hd__nand3_2 _32064_ (.A(_09716_),
    .B(_09717_),
    .C(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__a21o_1 _32065_ (.A1(_09488_),
    .A2(_09482_),
    .B1(_09487_),
    .X(_09721_));
 sky130_fd_sc_hd__buf_6 _32066_ (.A(_19595_),
    .X(_09722_));
 sky130_fd_sc_hd__buf_6 _32067_ (.A(_19599_),
    .X(_09723_));
 sky130_fd_sc_hd__a22oi_4 _32068_ (.A1(_09722_),
    .A2(_06020_),
    .B1(_09723_),
    .B2(_19924_),
    .Y(_09724_));
 sky130_fd_sc_hd__nor2_4 _32069_ (.A(_09714_),
    .B(_09715_),
    .Y(_09725_));
 sky130_fd_sc_hd__o21ai_2 _32070_ (.A1(_09724_),
    .A2(_09725_),
    .B1(_09718_),
    .Y(_09726_));
 sky130_fd_sc_hd__nand3_4 _32071_ (.A(_09720_),
    .B(_09721_),
    .C(_09726_),
    .Y(_09727_));
 sky130_fd_sc_hd__nand3_2 _32072_ (.A(_09716_),
    .B(_09717_),
    .C(_09718_),
    .Y(_09728_));
 sky130_fd_sc_hd__a21oi_2 _32073_ (.A1(_09488_),
    .A2(_09482_),
    .B1(_09487_),
    .Y(_09729_));
 sky130_fd_sc_hd__o21ai_2 _32074_ (.A1(_09724_),
    .A2(_09725_),
    .B1(_09719_),
    .Y(_09730_));
 sky130_fd_sc_hd__nand3_4 _32075_ (.A(_09728_),
    .B(_09729_),
    .C(_09730_),
    .Y(_09731_));
 sky130_fd_sc_hd__nand2_4 _32076_ (.A(_09727_),
    .B(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__a21oi_2 _32077_ (.A1(_09713_),
    .A2(_09732_),
    .B1(_09495_),
    .Y(_09733_));
 sky130_fd_sc_hd__nand3_4 _32078_ (.A(_09727_),
    .B(_09731_),
    .C(_09712_),
    .Y(_09734_));
 sky130_fd_sc_hd__nand2_1 _32079_ (.A(_09732_),
    .B(_09713_),
    .Y(_09735_));
 sky130_fd_sc_hd__a22oi_4 _32080_ (.A1(_09494_),
    .A2(_09491_),
    .B1(_09735_),
    .B2(_09734_),
    .Y(_09736_));
 sky130_fd_sc_hd__a21oi_4 _32081_ (.A1(_09733_),
    .A2(_09734_),
    .B1(_09736_),
    .Y(_09737_));
 sky130_fd_sc_hd__a21o_1 _32082_ (.A1(_09695_),
    .A2(_09701_),
    .B1(_09702_),
    .X(_09738_));
 sky130_fd_sc_hd__nand3_4 _32083_ (.A(_09695_),
    .B(_09702_),
    .C(_09701_),
    .Y(_09739_));
 sky130_fd_sc_hd__nand3_4 _32084_ (.A(_09738_),
    .B(_09739_),
    .C(_09705_),
    .Y(_09740_));
 sky130_fd_sc_hd__nand3_4 _32085_ (.A(_09707_),
    .B(_09737_),
    .C(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__and4_2 _32086_ (.A(_09735_),
    .B(_09494_),
    .C(_09491_),
    .D(_09734_),
    .X(_09742_));
 sky130_fd_sc_hd__nand3_2 _32087_ (.A(_09738_),
    .B(_09739_),
    .C(_09706_),
    .Y(_09743_));
 sky130_fd_sc_hd__o21ai_2 _32088_ (.A1(_09703_),
    .A2(_09704_),
    .B1(_09705_),
    .Y(_09744_));
 sky130_fd_sc_hd__o211ai_4 _32089_ (.A1(_09736_),
    .A2(_09742_),
    .B1(_09743_),
    .C1(_09744_),
    .Y(_09745_));
 sky130_fd_sc_hd__o2bb2ai_2 _32090_ (.A1_N(_09741_),
    .A2_N(_09745_),
    .B1(_09537_),
    .B2(_09545_),
    .Y(_09746_));
 sky130_fd_sc_hd__buf_2 _32091_ (.A(_09746_),
    .X(_09747_));
 sky130_fd_sc_hd__nand3b_4 _32092_ (.A_N(_09542_),
    .B(_09741_),
    .C(_09745_),
    .Y(_09748_));
 sky130_fd_sc_hd__nand2_1 _32093_ (.A(_09747_),
    .B(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__nand2_2 _32094_ (.A(_09672_),
    .B(_09749_),
    .Y(_09750_));
 sky130_fd_sc_hd__and3_2 _32095_ (.A(_09707_),
    .B(_09737_),
    .C(_09740_),
    .X(_09751_));
 sky130_fd_sc_hd__a21o_1 _32096_ (.A1(_09494_),
    .A2(_09491_),
    .B1(_09498_),
    .X(_09752_));
 sky130_fd_sc_hd__nor2_2 _32097_ (.A(_09752_),
    .B(_09531_),
    .Y(_09753_));
 sky130_fd_sc_hd__nand3_4 _32098_ (.A(_09745_),
    .B(_09753_),
    .C(_09540_),
    .Y(_09754_));
 sky130_fd_sc_hd__o2111ai_4 _32099_ (.A1(_09751_),
    .A2(_09754_),
    .B1(_09671_),
    .C1(_09747_),
    .D1(_09664_),
    .Y(_09755_));
 sky130_vsdinv _32100_ (.A(_09542_),
    .Y(_09756_));
 sky130_fd_sc_hd__nand2_1 _32101_ (.A(_09538_),
    .B(_09543_),
    .Y(_09757_));
 sky130_fd_sc_hd__o22ai_4 _32102_ (.A1(_09756_),
    .A2(_09757_),
    .B1(_09544_),
    .B2(_09562_),
    .Y(_09758_));
 sky130_fd_sc_hd__a21oi_4 _32103_ (.A1(_09750_),
    .A2(_09755_),
    .B1(_09758_),
    .Y(_09759_));
 sky130_vsdinv _32104_ (.A(_09664_),
    .Y(_09760_));
 sky130_fd_sc_hd__nand3_1 _32105_ (.A(_09747_),
    .B(_09748_),
    .C(_09671_),
    .Y(_09761_));
 sky130_fd_sc_hd__o211a_2 _32106_ (.A1(_09760_),
    .A2(_09761_),
    .B1(_09750_),
    .C1(_09758_),
    .X(_09762_));
 sky130_fd_sc_hd__a22oi_4 _32107_ (.A1(_05587_),
    .A2(_07705_),
    .B1(_05589_),
    .B2(_08336_),
    .Y(_09763_));
 sky130_vsdinv _32108_ (.A(_07686_),
    .Y(_09764_));
 sky130_fd_sc_hd__buf_4 _32109_ (.A(_09764_),
    .X(_09765_));
 sky130_fd_sc_hd__nand3_4 _32110_ (.A(_06492_),
    .B(_05447_),
    .C(_19868_),
    .Y(_09766_));
 sky130_fd_sc_hd__nor2_2 _32111_ (.A(_09765_),
    .B(_09766_),
    .Y(_09767_));
 sky130_fd_sc_hd__nand2_2 _32112_ (.A(_05835_),
    .B(_19862_),
    .Y(_09768_));
 sky130_fd_sc_hd__o21ai_2 _32113_ (.A1(_09763_),
    .A2(_09767_),
    .B1(_09768_),
    .Y(_09769_));
 sky130_fd_sc_hd__o21ai_2 _32114_ (.A1(_09449_),
    .A2(_09447_),
    .B1(_09453_),
    .Y(_09770_));
 sky130_vsdinv _32115_ (.A(_09768_),
    .Y(_09771_));
 sky130_fd_sc_hd__buf_4 _32116_ (.A(\pcpi_mul.rs1[21] ),
    .X(_09772_));
 sky130_fd_sc_hd__a22o_2 _32117_ (.A1(_06076_),
    .A2(_07701_),
    .B1(_06077_),
    .B2(_09772_),
    .X(_09773_));
 sky130_fd_sc_hd__o211ai_4 _32118_ (.A1(_09765_),
    .A2(_09766_),
    .B1(_09771_),
    .C1(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__nand3_4 _32119_ (.A(_09769_),
    .B(_09770_),
    .C(_09774_),
    .Y(_09775_));
 sky130_fd_sc_hd__o21ai_2 _32120_ (.A1(_09763_),
    .A2(_09767_),
    .B1(_09771_),
    .Y(_09776_));
 sky130_fd_sc_hd__a21oi_2 _32121_ (.A1(_09454_),
    .A2(_09450_),
    .B1(_09448_),
    .Y(_09777_));
 sky130_fd_sc_hd__o211ai_2 _32122_ (.A1(_09765_),
    .A2(_09766_),
    .B1(_09768_),
    .C1(_09773_),
    .Y(_09778_));
 sky130_fd_sc_hd__nand3_4 _32123_ (.A(_09776_),
    .B(_09777_),
    .C(_09778_),
    .Y(_09779_));
 sky130_fd_sc_hd__nor2_4 _32124_ (.A(_09314_),
    .B(_09311_),
    .Y(_09780_));
 sky130_fd_sc_hd__o2bb2ai_4 _32125_ (.A1_N(_09775_),
    .A2_N(_09779_),
    .B1(_09309_),
    .B2(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__nor2_4 _32126_ (.A(_09309_),
    .B(_09780_),
    .Y(_09782_));
 sky130_fd_sc_hd__nand3_4 _32127_ (.A(_09779_),
    .B(_09775_),
    .C(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__nand2_1 _32128_ (.A(_09445_),
    .B(_09456_),
    .Y(_09784_));
 sky130_fd_sc_hd__nand2_4 _32129_ (.A(_09784_),
    .B(_09444_),
    .Y(_09785_));
 sky130_fd_sc_hd__a21oi_4 _32130_ (.A1(_09781_),
    .A2(_09783_),
    .B1(_09785_),
    .Y(_09786_));
 sky130_vsdinv _32131_ (.A(_09775_),
    .Y(_09787_));
 sky130_fd_sc_hd__nand2_1 _32132_ (.A(_09779_),
    .B(_09782_),
    .Y(_09788_));
 sky130_fd_sc_hd__o211a_1 _32133_ (.A1(_09787_),
    .A2(_09788_),
    .B1(_09781_),
    .C1(_09785_),
    .X(_09789_));
 sky130_fd_sc_hd__nand2_1 _32134_ (.A(_09327_),
    .B(_09318_),
    .Y(_09790_));
 sky130_fd_sc_hd__o21ai_2 _32135_ (.A1(_09786_),
    .A2(_09789_),
    .B1(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__nand2_1 _32136_ (.A(_09328_),
    .B(_09336_),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_1 _32137_ (.A(_09792_),
    .B(_09330_),
    .Y(_09793_));
 sky130_fd_sc_hd__a21o_1 _32138_ (.A1(_09781_),
    .A2(_09783_),
    .B1(_09785_),
    .X(_09794_));
 sky130_fd_sc_hd__nand3_4 _32139_ (.A(_09785_),
    .B(_09781_),
    .C(_09783_),
    .Y(_09795_));
 sky130_fd_sc_hd__and2_2 _32140_ (.A(_09327_),
    .B(_09318_),
    .X(_09796_));
 sky130_fd_sc_hd__nand3_2 _32141_ (.A(_09794_),
    .B(_09795_),
    .C(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__nand3_4 _32142_ (.A(_09791_),
    .B(_09793_),
    .C(_09797_),
    .Y(_09798_));
 sky130_fd_sc_hd__o21ai_2 _32143_ (.A1(_09786_),
    .A2(_09789_),
    .B1(_09796_),
    .Y(_09799_));
 sky130_fd_sc_hd__a21oi_1 _32144_ (.A1(_09325_),
    .A2(_09327_),
    .B1(_09308_),
    .Y(_09800_));
 sky130_fd_sc_hd__o21ai_2 _32145_ (.A1(_09336_),
    .A2(_09800_),
    .B1(_09328_),
    .Y(_09801_));
 sky130_fd_sc_hd__nand3_2 _32146_ (.A(_09794_),
    .B(_09795_),
    .C(_09790_),
    .Y(_09802_));
 sky130_fd_sc_hd__nand3_4 _32147_ (.A(_09799_),
    .B(_09801_),
    .C(_09802_),
    .Y(_09803_));
 sky130_vsdinv _32148_ (.A(_19838_),
    .Y(_09804_));
 sky130_fd_sc_hd__buf_8 _32149_ (.A(_09804_),
    .X(_09805_));
 sky130_fd_sc_hd__buf_6 _32150_ (.A(_08487_),
    .X(_09806_));
 sky130_fd_sc_hd__nand3_4 _32151_ (.A(_05203_),
    .B(_05285_),
    .C(_08477_),
    .Y(_09807_));
 sky130_fd_sc_hd__a22o_1 _32152_ (.A1(_05772_),
    .A2(_08477_),
    .B1(_05562_),
    .B2(_09076_),
    .X(_09808_));
 sky130_fd_sc_hd__o21ai_2 _32153_ (.A1(_09806_),
    .A2(_09807_),
    .B1(_09808_),
    .Y(_09809_));
 sky130_fd_sc_hd__o21ai_4 _32154_ (.A1(_04839_),
    .A2(_09805_),
    .B1(_09809_),
    .Y(_09810_));
 sky130_fd_sc_hd__nor2_1 _32155_ (.A(_09806_),
    .B(_09807_),
    .Y(_09811_));
 sky130_fd_sc_hd__nor2_2 _32156_ (.A(_04838_),
    .B(_09804_),
    .Y(_09812_));
 sky130_fd_sc_hd__nand3b_4 _32157_ (.A_N(_09811_),
    .B(_09808_),
    .C(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__o21ai_4 _32158_ (.A1(_09351_),
    .A2(_09349_),
    .B1(_09348_),
    .Y(_09814_));
 sky130_fd_sc_hd__a21oi_4 _32159_ (.A1(_09810_),
    .A2(_09813_),
    .B1(_09814_),
    .Y(_09815_));
 sky130_fd_sc_hd__and3_1 _32160_ (.A(_09810_),
    .B(_09814_),
    .C(_09813_),
    .X(_09816_));
 sky130_fd_sc_hd__buf_6 _32161_ (.A(\pcpi_mul.rs1[27] ),
    .X(_09817_));
 sky130_fd_sc_hd__nand2_2 _32162_ (.A(_05233_),
    .B(_19848_),
    .Y(_09818_));
 sky130_fd_sc_hd__a21o_1 _32163_ (.A1(_05223_),
    .A2(_09817_),
    .B1(_09818_),
    .X(_09819_));
 sky130_fd_sc_hd__buf_4 _32164_ (.A(_19847_),
    .X(_09820_));
 sky130_fd_sc_hd__nand2_2 _32165_ (.A(_05227_),
    .B(_19843_),
    .Y(_09821_));
 sky130_fd_sc_hd__a21o_1 _32166_ (.A1(_06639_),
    .A2(_09820_),
    .B1(_09821_),
    .X(_09822_));
 sky130_fd_sc_hd__buf_6 _32167_ (.A(_09079_),
    .X(_09823_));
 sky130_fd_sc_hd__nand2_2 _32168_ (.A(_05157_),
    .B(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__a21oi_4 _32169_ (.A1(_09819_),
    .A2(_09822_),
    .B1(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__nand3_2 _32170_ (.A(_09819_),
    .B(_09822_),
    .C(_09824_),
    .Y(_09826_));
 sky130_vsdinv _32171_ (.A(_09826_),
    .Y(_09827_));
 sky130_fd_sc_hd__nor2_2 _32172_ (.A(_09825_),
    .B(_09827_),
    .Y(_09828_));
 sky130_fd_sc_hd__o21ai_2 _32173_ (.A1(_09815_),
    .A2(_09816_),
    .B1(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__a21boi_2 _32174_ (.A1(_09370_),
    .A2(_09376_),
    .B1_N(_09371_),
    .Y(_09830_));
 sky130_fd_sc_hd__a21o_1 _32175_ (.A1(_09810_),
    .A2(_09813_),
    .B1(_09814_),
    .X(_09831_));
 sky130_fd_sc_hd__a21o_1 _32176_ (.A1(_09819_),
    .A2(_09822_),
    .B1(_09824_),
    .X(_09832_));
 sky130_fd_sc_hd__nand2_2 _32177_ (.A(_09832_),
    .B(_09826_),
    .Y(_09833_));
 sky130_fd_sc_hd__nand3_4 _32178_ (.A(_09810_),
    .B(_09814_),
    .C(_09813_),
    .Y(_09834_));
 sky130_fd_sc_hd__nand3_2 _32179_ (.A(_09831_),
    .B(_09833_),
    .C(_09834_),
    .Y(_09835_));
 sky130_fd_sc_hd__nand3_4 _32180_ (.A(_09829_),
    .B(_09830_),
    .C(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__o22ai_4 _32181_ (.A1(_09825_),
    .A2(_09827_),
    .B1(_09815_),
    .B2(_09816_),
    .Y(_09837_));
 sky130_fd_sc_hd__nand3_2 _32182_ (.A(_09831_),
    .B(_09828_),
    .C(_09834_),
    .Y(_09838_));
 sky130_fd_sc_hd__o21ai_2 _32183_ (.A1(_09379_),
    .A2(_09357_),
    .B1(_09371_),
    .Y(_09839_));
 sky130_fd_sc_hd__nand3_4 _32184_ (.A(_09837_),
    .B(_09838_),
    .C(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__nor2_2 _32185_ (.A(_09360_),
    .B(_09363_),
    .Y(_09841_));
 sky130_fd_sc_hd__nor2_4 _32186_ (.A(_09841_),
    .B(_09367_),
    .Y(_09842_));
 sky130_vsdinv _32187_ (.A(_09842_),
    .Y(_09843_));
 sky130_fd_sc_hd__and3_1 _32188_ (.A(_09836_),
    .B(_09840_),
    .C(_09843_),
    .X(_09844_));
 sky130_fd_sc_hd__nand2_1 _32189_ (.A(_09836_),
    .B(_09840_),
    .Y(_09845_));
 sky130_fd_sc_hd__and2_1 _32190_ (.A(_09845_),
    .B(_09842_),
    .X(_09846_));
 sky130_fd_sc_hd__o2bb2ai_4 _32191_ (.A1_N(_09798_),
    .A2_N(_09803_),
    .B1(_09844_),
    .B2(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__nand2_2 _32192_ (.A(_09549_),
    .B(_09472_),
    .Y(_09848_));
 sky130_fd_sc_hd__nand2_1 _32193_ (.A(_09845_),
    .B(_09843_),
    .Y(_09849_));
 sky130_fd_sc_hd__nand3_1 _32194_ (.A(_09836_),
    .B(_09840_),
    .C(_09842_),
    .Y(_09850_));
 sky130_fd_sc_hd__nand2_2 _32195_ (.A(_09849_),
    .B(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__nand3_4 _32196_ (.A(_09851_),
    .B(_09803_),
    .C(_09798_),
    .Y(_09852_));
 sky130_fd_sc_hd__nand3_4 _32197_ (.A(_09847_),
    .B(_09848_),
    .C(_09852_),
    .Y(_09853_));
 sky130_vsdinv _32198_ (.A(_09344_),
    .Y(_09854_));
 sky130_fd_sc_hd__a21oi_4 _32199_ (.A1(_09391_),
    .A2(_09338_),
    .B1(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__a21oi_4 _32200_ (.A1(_09847_),
    .A2(_09852_),
    .B1(_09848_),
    .Y(_09856_));
 sky130_fd_sc_hd__nor2_2 _32201_ (.A(_09855_),
    .B(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__a21oi_2 _32202_ (.A1(_09803_),
    .A2(_09798_),
    .B1(_09851_),
    .Y(_09858_));
 sky130_fd_sc_hd__a21oi_1 _32203_ (.A1(_09836_),
    .A2(_09840_),
    .B1(_09842_),
    .Y(_09859_));
 sky130_fd_sc_hd__and3_1 _32204_ (.A(_09836_),
    .B(_09840_),
    .C(_09842_),
    .X(_09860_));
 sky130_fd_sc_hd__o211a_1 _32205_ (.A1(_09859_),
    .A2(_09860_),
    .B1(_09798_),
    .C1(_09803_),
    .X(_09861_));
 sky130_fd_sc_hd__o21bai_4 _32206_ (.A1(_09858_),
    .A2(_09861_),
    .B1_N(_09848_),
    .Y(_09862_));
 sky130_fd_sc_hd__a21o_2 _32207_ (.A1(_09391_),
    .A2(_09338_),
    .B1(_09854_),
    .X(_09863_));
 sky130_fd_sc_hd__a21oi_4 _32208_ (.A1(_09862_),
    .A2(_09853_),
    .B1(_09863_),
    .Y(_09864_));
 sky130_fd_sc_hd__a21oi_1 _32209_ (.A1(_09853_),
    .A2(_09857_),
    .B1(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__o21ai_2 _32210_ (.A1(_09759_),
    .A2(_09762_),
    .B1(_09865_),
    .Y(_09866_));
 sky130_fd_sc_hd__a21o_1 _32211_ (.A1(_09396_),
    .A2(_09400_),
    .B1(_09402_),
    .X(_09867_));
 sky130_fd_sc_hd__nand3_4 _32212_ (.A(_09396_),
    .B(_09400_),
    .C(_09402_),
    .Y(_09868_));
 sky130_fd_sc_hd__a21oi_2 _32213_ (.A1(_09559_),
    .A2(_09563_),
    .B1(_09561_),
    .Y(_09869_));
 sky130_fd_sc_hd__a31oi_4 _32214_ (.A1(_09564_),
    .A2(_09867_),
    .A3(_09868_),
    .B1(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__o211a_4 _32215_ (.A1(_09548_),
    .A2(_09557_),
    .B1(_09852_),
    .C1(_09847_),
    .X(_09871_));
 sky130_fd_sc_hd__o21ai_4 _32216_ (.A1(_09856_),
    .A2(_09871_),
    .B1(_09855_),
    .Y(_09872_));
 sky130_fd_sc_hd__nand3_4 _32217_ (.A(_09862_),
    .B(_09853_),
    .C(_09863_),
    .Y(_09873_));
 sky130_fd_sc_hd__nand2_2 _32218_ (.A(_09872_),
    .B(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__a22oi_4 _32219_ (.A1(_09747_),
    .A2(_09748_),
    .B1(_09664_),
    .B2(_09671_),
    .Y(_09875_));
 sky130_fd_sc_hd__o2111a_1 _32220_ (.A1(_09751_),
    .A2(_09754_),
    .B1(_09671_),
    .C1(_09747_),
    .D1(_09664_),
    .X(_09876_));
 sky130_fd_sc_hd__a21oi_4 _32221_ (.A1(_09558_),
    .A2(_09553_),
    .B1(_09546_),
    .Y(_09877_));
 sky130_fd_sc_hd__o21ai_4 _32222_ (.A1(_09875_),
    .A2(_09876_),
    .B1(_09877_),
    .Y(_09878_));
 sky130_fd_sc_hd__nand3_4 _32223_ (.A(_09758_),
    .B(_09750_),
    .C(_09755_),
    .Y(_09879_));
 sky130_fd_sc_hd__nand3_4 _32224_ (.A(_09874_),
    .B(_09878_),
    .C(_09879_),
    .Y(_09880_));
 sky130_fd_sc_hd__nand3_4 _32225_ (.A(_09866_),
    .B(_09870_),
    .C(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__and3_1 _32226_ (.A(_09862_),
    .B(_09853_),
    .C(_09863_),
    .X(_09882_));
 sky130_fd_sc_hd__o22ai_4 _32227_ (.A1(_09864_),
    .A2(_09882_),
    .B1(_09759_),
    .B2(_09762_),
    .Y(_09883_));
 sky130_fd_sc_hd__nand2_2 _32228_ (.A(_09862_),
    .B(_09863_),
    .Y(_09884_));
 sky130_fd_sc_hd__o2111ai_4 _32229_ (.A1(_09871_),
    .A2(_09884_),
    .B1(_09872_),
    .C1(_09879_),
    .D1(_09878_),
    .Y(_09885_));
 sky130_fd_sc_hd__nand3_1 _32230_ (.A(_09564_),
    .B(_09867_),
    .C(_09868_),
    .Y(_09886_));
 sky130_fd_sc_hd__nand2_2 _32231_ (.A(_09886_),
    .B(_09555_),
    .Y(_09887_));
 sky130_fd_sc_hd__nand3_4 _32232_ (.A(_09883_),
    .B(_09885_),
    .C(_09887_),
    .Y(_09888_));
 sky130_vsdinv _32233_ (.A(_09388_),
    .Y(_09889_));
 sky130_fd_sc_hd__nand2_4 _32234_ (.A(_09889_),
    .B(_09383_),
    .Y(_09890_));
 sky130_fd_sc_hd__nand2_1 _32235_ (.A(_09396_),
    .B(_09402_),
    .Y(_09891_));
 sky130_fd_sc_hd__nand2_4 _32236_ (.A(_09891_),
    .B(_09400_),
    .Y(_09892_));
 sky130_fd_sc_hd__nor2_8 _32237_ (.A(_09890_),
    .B(_09892_),
    .Y(_09893_));
 sky130_vsdinv _32238_ (.A(_09890_),
    .Y(_09894_));
 sky130_vsdinv _32239_ (.A(_09892_),
    .Y(_09895_));
 sky130_fd_sc_hd__nor2_8 _32240_ (.A(_09894_),
    .B(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__nor2_8 _32241_ (.A(_09893_),
    .B(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__a21oi_4 _32242_ (.A1(_09881_),
    .A2(_09888_),
    .B1(_09897_),
    .Y(_09898_));
 sky130_fd_sc_hd__a21oi_4 _32243_ (.A1(_09570_),
    .A2(_09571_),
    .B1(_09569_),
    .Y(_09899_));
 sky130_fd_sc_hd__nand3_2 _32244_ (.A(_09881_),
    .B(_09888_),
    .C(_09897_),
    .Y(_09900_));
 sky130_fd_sc_hd__o21ai_4 _32245_ (.A1(_09899_),
    .A2(_09580_),
    .B1(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__nor2_1 _32246_ (.A(_09890_),
    .B(_09895_),
    .Y(_09902_));
 sky130_fd_sc_hd__nor2_1 _32247_ (.A(_09894_),
    .B(_09892_),
    .Y(_09903_));
 sky130_fd_sc_hd__o2bb2ai_2 _32248_ (.A1_N(_09888_),
    .A2_N(_09881_),
    .B1(_09902_),
    .B2(_09903_),
    .Y(_09904_));
 sky130_fd_sc_hd__a21oi_2 _32249_ (.A1(_09572_),
    .A2(_09585_),
    .B1(_09899_),
    .Y(_09905_));
 sky130_fd_sc_hd__o211ai_4 _32250_ (.A1(_09896_),
    .A2(_09893_),
    .B1(_09888_),
    .C1(_09881_),
    .Y(_09906_));
 sky130_fd_sc_hd__nand3_4 _32251_ (.A(_09904_),
    .B(_09905_),
    .C(_09906_),
    .Y(_09907_));
 sky130_fd_sc_hd__o211ai_4 _32252_ (.A1(_09898_),
    .A2(_09901_),
    .B1(_09575_),
    .C1(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__o21ai_2 _32253_ (.A1(_09898_),
    .A2(_09901_),
    .B1(_09907_),
    .Y(_09909_));
 sky130_vsdinv _32254_ (.A(_09575_),
    .Y(_09910_));
 sky130_fd_sc_hd__nand2_2 _32255_ (.A(_09909_),
    .B(_09910_),
    .Y(_09911_));
 sky130_fd_sc_hd__a21oi_4 _32256_ (.A1(_09586_),
    .A2(_09584_),
    .B1(_09583_),
    .Y(_09912_));
 sky130_vsdinv _32257_ (.A(_09016_),
    .Y(_09913_));
 sky130_fd_sc_hd__a31oi_4 _32258_ (.A1(_09583_),
    .A2(_09586_),
    .A3(_09584_),
    .B1(_09913_),
    .Y(_09914_));
 sky130_fd_sc_hd__o2bb2ai_2 _32259_ (.A1_N(_09908_),
    .A2_N(_09911_),
    .B1(_09912_),
    .B2(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__a21oi_4 _32260_ (.A1(_09587_),
    .A2(_09016_),
    .B1(_09912_),
    .Y(_09916_));
 sky130_fd_sc_hd__nand3_4 _32261_ (.A(_09916_),
    .B(_09911_),
    .C(_09908_),
    .Y(_09917_));
 sky130_fd_sc_hd__nand2_1 _32262_ (.A(_09915_),
    .B(_09917_),
    .Y(_09918_));
 sky130_fd_sc_hd__nand3_4 _32263_ (.A(_09302_),
    .B(_09300_),
    .C(_09596_),
    .Y(_09919_));
 sky130_vsdinv _32264_ (.A(_09919_),
    .Y(_09920_));
 sky130_vsdinv _32265_ (.A(_09592_),
    .Y(_09921_));
 sky130_fd_sc_hd__a21oi_2 _32266_ (.A1(_09921_),
    .A2(_09299_),
    .B1(_09595_),
    .Y(_09922_));
 sky130_fd_sc_hd__nand3_2 _32267_ (.A(_09300_),
    .B(_09596_),
    .C(_09303_),
    .Y(_09923_));
 sky130_fd_sc_hd__nand2_4 _32268_ (.A(_09922_),
    .B(_09923_),
    .Y(_09924_));
 sky130_fd_sc_hd__a21oi_4 _32269_ (.A1(_09301_),
    .A2(_09920_),
    .B1(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__xor2_2 _32270_ (.A(_09918_),
    .B(_09925_),
    .X(_02647_));
 sky130_fd_sc_hd__a2bb2oi_4 _32271_ (.A1_N(_09898_),
    .A2_N(_09901_),
    .B1(_09910_),
    .B2(_09907_),
    .Y(_09926_));
 sky130_fd_sc_hd__and2_1 _32272_ (.A(_09668_),
    .B(_09467_),
    .X(_09927_));
 sky130_fd_sc_hd__nand2_2 _32273_ (.A(_09927_),
    .B(_09667_),
    .Y(_09928_));
 sky130_fd_sc_hd__buf_6 _32274_ (.A(_09806_),
    .X(_09929_));
 sky130_fd_sc_hd__nand2_2 _32275_ (.A(_05280_),
    .B(_09076_),
    .Y(_09930_));
 sky130_fd_sc_hd__nand2_2 _32276_ (.A(_05366_),
    .B(_09079_),
    .Y(_09931_));
 sky130_fd_sc_hd__or2_2 _32277_ (.A(_09930_),
    .B(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__clkbuf_4 _32278_ (.A(\pcpi_mul.rs1[29] ),
    .X(_09933_));
 sky130_fd_sc_hd__nand2_2 _32279_ (.A(_05171_),
    .B(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__nand2_2 _32280_ (.A(_09930_),
    .B(_09931_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand3_2 _32281_ (.A(_09932_),
    .B(_09934_),
    .C(_09935_),
    .Y(_09936_));
 sky130_fd_sc_hd__nor2_4 _32282_ (.A(_09930_),
    .B(_09931_),
    .Y(_09937_));
 sky130_fd_sc_hd__and2_1 _32283_ (.A(_09930_),
    .B(_09931_),
    .X(_09938_));
 sky130_vsdinv _32284_ (.A(_09934_),
    .Y(_09939_));
 sky130_fd_sc_hd__o21ai_2 _32285_ (.A1(_09937_),
    .A2(_09938_),
    .B1(_09939_),
    .Y(_09940_));
 sky130_fd_sc_hd__o2111ai_4 _32286_ (.A1(_09929_),
    .A2(_09807_),
    .B1(_09813_),
    .C1(_09936_),
    .D1(_09940_),
    .Y(_09941_));
 sky130_fd_sc_hd__a21o_1 _32287_ (.A1(_09812_),
    .A2(_09808_),
    .B1(_09811_),
    .X(_09942_));
 sky130_fd_sc_hd__o21ai_2 _32288_ (.A1(_09937_),
    .A2(_09938_),
    .B1(_09934_),
    .Y(_09943_));
 sky130_fd_sc_hd__nand3_2 _32289_ (.A(_09932_),
    .B(_09939_),
    .C(_09935_),
    .Y(_09944_));
 sky130_fd_sc_hd__nand3_4 _32290_ (.A(_09942_),
    .B(_09943_),
    .C(_09944_),
    .Y(_09945_));
 sky130_fd_sc_hd__buf_4 _32291_ (.A(\pcpi_mul.rs1[28] ),
    .X(_09946_));
 sky130_fd_sc_hd__clkbuf_4 _32292_ (.A(\pcpi_mul.rs1[27] ),
    .X(_09947_));
 sky130_fd_sc_hd__nand2_2 _32293_ (.A(_05266_),
    .B(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__a21o_1 _32294_ (.A1(_05239_),
    .A2(_09946_),
    .B1(_09948_),
    .X(_09949_));
 sky130_fd_sc_hd__buf_4 _32295_ (.A(_09947_),
    .X(_09950_));
 sky130_fd_sc_hd__nand2_2 _32296_ (.A(_05152_),
    .B(_19838_),
    .Y(_09951_));
 sky130_fd_sc_hd__a21o_1 _32297_ (.A1(_19679_),
    .A2(_09950_),
    .B1(_09951_),
    .X(_09952_));
 sky130_fd_sc_hd__nand2_2 _32298_ (.A(_05670_),
    .B(_09820_),
    .Y(_09953_));
 sky130_fd_sc_hd__a21oi_4 _32299_ (.A1(_09949_),
    .A2(_09952_),
    .B1(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__and3_2 _32300_ (.A(_09949_),
    .B(_09952_),
    .C(_09953_),
    .X(_09955_));
 sky130_fd_sc_hd__nor2_8 _32301_ (.A(_09954_),
    .B(_09955_),
    .Y(_09956_));
 sky130_fd_sc_hd__a21o_1 _32302_ (.A1(_09941_),
    .A2(_09945_),
    .B1(_09956_),
    .X(_09957_));
 sky130_fd_sc_hd__nand3_4 _32303_ (.A(_09956_),
    .B(_09941_),
    .C(_09945_),
    .Y(_09958_));
 sky130_fd_sc_hd__o21ai_4 _32304_ (.A1(_09833_),
    .A2(_09815_),
    .B1(_09834_),
    .Y(_09959_));
 sky130_fd_sc_hd__a21o_1 _32305_ (.A1(_09957_),
    .A2(_09958_),
    .B1(_09959_),
    .X(_09960_));
 sky130_fd_sc_hd__nand3_4 _32306_ (.A(_09957_),
    .B(_09959_),
    .C(_09958_),
    .Y(_09961_));
 sky130_fd_sc_hd__o21ai_4 _32307_ (.A1(_09818_),
    .A2(_09821_),
    .B1(_09832_),
    .Y(_09962_));
 sky130_fd_sc_hd__a21oi_2 _32308_ (.A1(_09960_),
    .A2(_09961_),
    .B1(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__and3_1 _32309_ (.A(_09957_),
    .B(_09959_),
    .C(_09958_),
    .X(_09964_));
 sky130_fd_sc_hd__nand2_2 _32310_ (.A(_09960_),
    .B(_09962_),
    .Y(_09965_));
 sky130_fd_sc_hd__nor2_2 _32311_ (.A(_09964_),
    .B(_09965_),
    .Y(_09966_));
 sky130_vsdinv _32312_ (.A(_09779_),
    .Y(_09967_));
 sky130_fd_sc_hd__nor2_2 _32313_ (.A(_09782_),
    .B(_09787_),
    .Y(_09968_));
 sky130_fd_sc_hd__a22oi_4 _32314_ (.A1(_19662_),
    .A2(_08333_),
    .B1(_06504_),
    .B2(_08337_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand3_4 _32315_ (.A(_05591_),
    .B(_19664_),
    .C(_19865_),
    .Y(_09970_));
 sky130_fd_sc_hd__nor2_2 _32316_ (.A(_08043_),
    .B(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__buf_4 _32317_ (.A(\pcpi_mul.rs1[23] ),
    .X(_09972_));
 sky130_fd_sc_hd__nand2_2 _32318_ (.A(_05443_),
    .B(_09972_),
    .Y(_09973_));
 sky130_vsdinv _32319_ (.A(_09973_),
    .Y(_09974_));
 sky130_fd_sc_hd__o21ai_2 _32320_ (.A1(_09969_),
    .A2(_09971_),
    .B1(_09974_),
    .Y(_09975_));
 sky130_fd_sc_hd__a21oi_2 _32321_ (.A1(_09609_),
    .A2(_09604_),
    .B1(_09602_),
    .Y(_09976_));
 sky130_fd_sc_hd__a22o_2 _32322_ (.A1(_05451_),
    .A2(_08056_),
    .B1(_05833_),
    .B2(_19862_),
    .X(_09977_));
 sky130_fd_sc_hd__o211ai_2 _32323_ (.A1(_08043_),
    .A2(_09970_),
    .B1(_09973_),
    .C1(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__nand3_4 _32324_ (.A(_09975_),
    .B(_09976_),
    .C(_09978_),
    .Y(_09979_));
 sky130_fd_sc_hd__o21ai_2 _32325_ (.A1(_09969_),
    .A2(_09971_),
    .B1(_09973_),
    .Y(_09980_));
 sky130_fd_sc_hd__o211ai_4 _32326_ (.A1(_08043_),
    .A2(_09970_),
    .B1(_09974_),
    .C1(_09977_),
    .Y(_09981_));
 sky130_fd_sc_hd__o21ai_2 _32327_ (.A1(_09603_),
    .A2(_09601_),
    .B1(_09608_),
    .Y(_09982_));
 sky130_fd_sc_hd__nand3_4 _32328_ (.A(_09980_),
    .B(_09981_),
    .C(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__a21o_2 _32329_ (.A1(_09773_),
    .A2(_09771_),
    .B1(_09767_),
    .X(_09984_));
 sky130_fd_sc_hd__a21o_2 _32330_ (.A1(_09979_),
    .A2(_09983_),
    .B1(_09984_),
    .X(_09985_));
 sky130_fd_sc_hd__nand3_4 _32331_ (.A(_09979_),
    .B(_09983_),
    .C(_09984_),
    .Y(_09986_));
 sky130_fd_sc_hd__nand2_1 _32332_ (.A(_09624_),
    .B(_09611_),
    .Y(_09987_));
 sky130_fd_sc_hd__nand2_4 _32333_ (.A(_09987_),
    .B(_09621_),
    .Y(_09988_));
 sky130_fd_sc_hd__a21oi_4 _32334_ (.A1(_09985_),
    .A2(_09986_),
    .B1(_09988_),
    .Y(_09989_));
 sky130_fd_sc_hd__and3_1 _32335_ (.A(_09980_),
    .B(_09982_),
    .C(_09981_),
    .X(_09990_));
 sky130_fd_sc_hd__nand2_1 _32336_ (.A(_09979_),
    .B(_09984_),
    .Y(_09991_));
 sky130_fd_sc_hd__o211a_1 _32337_ (.A1(_09990_),
    .A2(_09991_),
    .B1(_09985_),
    .C1(_09988_),
    .X(_09992_));
 sky130_fd_sc_hd__o22ai_4 _32338_ (.A1(_09967_),
    .A2(_09968_),
    .B1(_09989_),
    .B2(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__a21oi_2 _32339_ (.A1(_09979_),
    .A2(_09983_),
    .B1(_09984_),
    .Y(_09994_));
 sky130_vsdinv _32340_ (.A(_09986_),
    .Y(_09995_));
 sky130_fd_sc_hd__o21bai_4 _32341_ (.A1(_09994_),
    .A2(_09995_),
    .B1_N(_09988_),
    .Y(_09996_));
 sky130_fd_sc_hd__nand3_4 _32342_ (.A(_09988_),
    .B(_09985_),
    .C(_09986_),
    .Y(_09997_));
 sky130_fd_sc_hd__nand2_2 _32343_ (.A(_09788_),
    .B(_09775_),
    .Y(_09998_));
 sky130_fd_sc_hd__nand3_4 _32344_ (.A(_09996_),
    .B(_09997_),
    .C(_09998_),
    .Y(_09999_));
 sky130_fd_sc_hd__o21ai_4 _32345_ (.A1(_09796_),
    .A2(_09786_),
    .B1(_09795_),
    .Y(_10000_));
 sky130_fd_sc_hd__a21oi_2 _32346_ (.A1(_09993_),
    .A2(_09999_),
    .B1(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__nor2_1 _32347_ (.A(_09796_),
    .B(_09786_),
    .Y(_10002_));
 sky130_fd_sc_hd__o211a_2 _32348_ (.A1(_09789_),
    .A2(_10002_),
    .B1(_09999_),
    .C1(_09993_),
    .X(_10003_));
 sky130_fd_sc_hd__o22ai_4 _32349_ (.A1(_09963_),
    .A2(_09966_),
    .B1(_10001_),
    .B2(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__a21o_1 _32350_ (.A1(_09993_),
    .A2(_09999_),
    .B1(_10000_),
    .X(_10005_));
 sky130_fd_sc_hd__a21oi_1 _32351_ (.A1(_09957_),
    .A2(_09958_),
    .B1(_09959_),
    .Y(_10006_));
 sky130_fd_sc_hd__o21ai_1 _32352_ (.A1(_10006_),
    .A2(_09964_),
    .B1(_09962_),
    .Y(_10007_));
 sky130_fd_sc_hd__nand3b_1 _32353_ (.A_N(_09962_),
    .B(_09960_),
    .C(_09961_),
    .Y(_10008_));
 sky130_fd_sc_hd__nand2_2 _32354_ (.A(_10007_),
    .B(_10008_),
    .Y(_10009_));
 sky130_fd_sc_hd__nand3_4 _32355_ (.A(_09993_),
    .B(_10000_),
    .C(_09999_),
    .Y(_10010_));
 sky130_fd_sc_hd__nand3_4 _32356_ (.A(_10005_),
    .B(_10009_),
    .C(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__a22oi_4 _32357_ (.A1(_09666_),
    .A2(_09928_),
    .B1(_10004_),
    .B2(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__nor2_4 _32358_ (.A(_09927_),
    .B(_09660_),
    .Y(_10013_));
 sky130_fd_sc_hd__o211a_4 _32359_ (.A1(_09662_),
    .A2(_10013_),
    .B1(_10011_),
    .C1(_10004_),
    .X(_10014_));
 sky130_vsdinv _32360_ (.A(_09803_),
    .Y(_10015_));
 sky130_fd_sc_hd__a21o_2 _32361_ (.A1(_09798_),
    .A2(_09851_),
    .B1(_10015_),
    .X(_10016_));
 sky130_vsdinv _32362_ (.A(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__o21ai_4 _32363_ (.A1(_10012_),
    .A2(_10014_),
    .B1(_10017_),
    .Y(_10018_));
 sky130_vsdinv _32364_ (.A(_09928_),
    .Y(_10019_));
 sky130_fd_sc_hd__o2bb2ai_2 _32365_ (.A1_N(_10011_),
    .A2_N(_10004_),
    .B1(_09660_),
    .B2(_10019_),
    .Y(_10020_));
 sky130_fd_sc_hd__o211ai_4 _32366_ (.A1(_09662_),
    .A2(_10013_),
    .B1(_10011_),
    .C1(_10004_),
    .Y(_10021_));
 sky130_fd_sc_hd__nand3_4 _32367_ (.A(_10020_),
    .B(_10021_),
    .C(_10016_),
    .Y(_10022_));
 sky130_fd_sc_hd__nand2_1 _32368_ (.A(_10018_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__nand3_1 _32369_ (.A(_09664_),
    .B(_09670_),
    .C(_09747_),
    .Y(_10024_));
 sky130_fd_sc_hd__nand2_2 _32370_ (.A(_10024_),
    .B(_09748_),
    .Y(_10025_));
 sky130_fd_sc_hd__nand3_4 _32371_ (.A(\pcpi_mul.rs2[26] ),
    .B(\pcpi_mul.rs2[25] ),
    .C(_05172_),
    .Y(_10026_));
 sky130_fd_sc_hd__nor2_4 _32372_ (.A(_05154_),
    .B(_10026_),
    .Y(_10027_));
 sky130_fd_sc_hd__nand2_2 _32373_ (.A(\pcpi_mul.rs2[24] ),
    .B(_19916_),
    .Y(_10028_));
 sky130_fd_sc_hd__a22o_2 _32374_ (.A1(_09229_),
    .A2(_05695_),
    .B1(_19599_),
    .B2(_07008_),
    .X(_10029_));
 sky130_fd_sc_hd__nand3b_4 _32375_ (.A_N(_10027_),
    .B(_10028_),
    .C(_10029_),
    .Y(_10030_));
 sky130_vsdinv _32376_ (.A(_09710_),
    .Y(_10031_));
 sky130_fd_sc_hd__a22oi_4 _32377_ (.A1(_19596_),
    .A2(_05146_),
    .B1(_09227_),
    .B2(_05224_),
    .Y(_10032_));
 sky130_vsdinv _32378_ (.A(_10028_),
    .Y(_10033_));
 sky130_fd_sc_hd__o21ai_2 _32379_ (.A1(_10032_),
    .A2(_10027_),
    .B1(_10033_),
    .Y(_10034_));
 sky130_fd_sc_hd__nand3_2 _32380_ (.A(_10030_),
    .B(_10031_),
    .C(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__nand3b_2 _32381_ (.A_N(_10027_),
    .B(_10033_),
    .C(_10029_),
    .Y(_10036_));
 sky130_fd_sc_hd__o21ai_2 _32382_ (.A1(_10032_),
    .A2(_10027_),
    .B1(_10028_),
    .Y(_10037_));
 sky130_fd_sc_hd__nand3_4 _32383_ (.A(_10036_),
    .B(_09710_),
    .C(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__nand2_1 _32384_ (.A(_10035_),
    .B(_10038_),
    .Y(_10039_));
 sky130_fd_sc_hd__a21oi_4 _32385_ (.A1(_09719_),
    .A2(_09717_),
    .B1(_09725_),
    .Y(_10040_));
 sky130_fd_sc_hd__nand2_4 _32386_ (.A(_10039_),
    .B(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__a31oi_4 _32387_ (.A1(_10030_),
    .A2(_10034_),
    .A3(_10031_),
    .B1(_10040_),
    .Y(_10042_));
 sky130_fd_sc_hd__nand2_4 _32388_ (.A(_10042_),
    .B(_10038_),
    .Y(_10043_));
 sky130_vsdinv _32389_ (.A(\pcpi_mul.rs2[27] ),
    .Y(_10044_));
 sky130_fd_sc_hd__nor2_8 _32390_ (.A(_10044_),
    .B(_05150_),
    .Y(_10045_));
 sky130_fd_sc_hd__buf_6 _32391_ (.A(\pcpi_mul.rs2[28] ),
    .X(_10046_));
 sky130_fd_sc_hd__nand2_2 _32392_ (.A(_10046_),
    .B(_05441_),
    .Y(_10047_));
 sky130_fd_sc_hd__nand2_2 _32393_ (.A(_19582_),
    .B(_05204_),
    .Y(_10048_));
 sky130_fd_sc_hd__nor2_4 _32394_ (.A(_10047_),
    .B(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__and2_1 _32395_ (.A(_10047_),
    .B(_10048_),
    .X(_10050_));
 sky130_fd_sc_hd__nor2_4 _32396_ (.A(_10049_),
    .B(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__xor2_4 _32397_ (.A(_10045_),
    .B(_10051_),
    .X(_10052_));
 sky130_fd_sc_hd__a21oi_4 _32398_ (.A1(_10041_),
    .A2(_10043_),
    .B1(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__and3_4 _32399_ (.A(_10041_),
    .B(_10043_),
    .C(_10052_),
    .X(_10054_));
 sky130_fd_sc_hd__o22ai_4 _32400_ (.A1(_09713_),
    .A2(_09732_),
    .B1(_10053_),
    .B2(_10054_),
    .Y(_10055_));
 sky130_fd_sc_hd__nand2_2 _32401_ (.A(_10041_),
    .B(_10043_),
    .Y(_10056_));
 sky130_vsdinv _32402_ (.A(_10052_),
    .Y(_10057_));
 sky130_fd_sc_hd__nand2_4 _32403_ (.A(_10056_),
    .B(_10057_),
    .Y(_10058_));
 sky130_vsdinv _32404_ (.A(_09734_),
    .Y(_10059_));
 sky130_fd_sc_hd__nand3_4 _32405_ (.A(_10041_),
    .B(_10052_),
    .C(_10043_),
    .Y(_10060_));
 sky130_fd_sc_hd__nand3_4 _32406_ (.A(_10058_),
    .B(_10059_),
    .C(_10060_),
    .Y(_10061_));
 sky130_fd_sc_hd__nand2_2 _32407_ (.A(_10055_),
    .B(_10061_),
    .Y(_10062_));
 sky130_vsdinv _32408_ (.A(_09687_),
    .Y(_10063_));
 sky130_fd_sc_hd__and3_1 _32409_ (.A(_09683_),
    .B(_09698_),
    .C(_09699_),
    .X(_10064_));
 sky130_fd_sc_hd__o22ai_4 _32410_ (.A1(_05278_),
    .A2(_09674_),
    .B1(_09676_),
    .B2(_09673_),
    .Y(_10065_));
 sky130_fd_sc_hd__buf_4 _32411_ (.A(_09516_),
    .X(_10066_));
 sky130_fd_sc_hd__a22oi_4 _32412_ (.A1(_08549_),
    .A2(_05637_),
    .B1(_10066_),
    .B2(_08198_),
    .Y(_10067_));
 sky130_fd_sc_hd__nand3_4 _32413_ (.A(_08539_),
    .B(_09516_),
    .C(_05483_),
    .Y(_10068_));
 sky130_fd_sc_hd__nor2_4 _32414_ (.A(_08197_),
    .B(_10068_),
    .Y(_10069_));
 sky130_fd_sc_hd__nand2_4 _32415_ (.A(_08545_),
    .B(_19906_),
    .Y(_10070_));
 sky130_vsdinv _32416_ (.A(_10070_),
    .Y(_10071_));
 sky130_fd_sc_hd__o21ai_2 _32417_ (.A1(_10067_),
    .A2(_10069_),
    .B1(_10071_),
    .Y(_10072_));
 sky130_fd_sc_hd__buf_2 _32418_ (.A(_19606_),
    .X(_10073_));
 sky130_fd_sc_hd__a22o_2 _32419_ (.A1(_10073_),
    .A2(_05291_),
    .B1(_09680_),
    .B2(_08198_),
    .X(_10074_));
 sky130_fd_sc_hd__o211ai_4 _32420_ (.A1(_08197_),
    .A2(_10068_),
    .B1(_10070_),
    .C1(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__nand3b_4 _32421_ (.A_N(_10065_),
    .B(_10072_),
    .C(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__o21ai_2 _32422_ (.A1(_10067_),
    .A2(_10069_),
    .B1(_10070_),
    .Y(_10077_));
 sky130_fd_sc_hd__o211ai_4 _32423_ (.A1(_08197_),
    .A2(_10068_),
    .B1(_10071_),
    .C1(_10074_),
    .Y(_10078_));
 sky130_fd_sc_hd__nand3_4 _32424_ (.A(_10077_),
    .B(_10065_),
    .C(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__a22oi_2 _32425_ (.A1(_07486_),
    .A2(_05673_),
    .B1(_08172_),
    .B2(_06441_),
    .Y(_10080_));
 sky130_fd_sc_hd__nand2_2 _32426_ (.A(_07822_),
    .B(_05558_),
    .Y(_10081_));
 sky130_fd_sc_hd__nand2_2 _32427_ (.A(_07824_),
    .B(_06259_),
    .Y(_10082_));
 sky130_fd_sc_hd__nor2_4 _32428_ (.A(_10081_),
    .B(_10082_),
    .Y(_10083_));
 sky130_fd_sc_hd__nor2_1 _32429_ (.A(_10080_),
    .B(_10083_),
    .Y(_10084_));
 sky130_fd_sc_hd__o21ai_1 _32430_ (.A1(_07042_),
    .A2(_05788_),
    .B1(_10084_),
    .Y(_10085_));
 sky130_fd_sc_hd__nor2_1 _32431_ (.A(_07041_),
    .B(_07102_),
    .Y(_10086_));
 sky130_fd_sc_hd__o21ai_1 _32432_ (.A1(_10080_),
    .A2(_10083_),
    .B1(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__nand2_2 _32433_ (.A(_10085_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__a21o_2 _32434_ (.A1(_10076_),
    .A2(_10079_),
    .B1(_10088_),
    .X(_10089_));
 sky130_fd_sc_hd__nand3_4 _32435_ (.A(_10088_),
    .B(_10079_),
    .C(_10076_),
    .Y(_10090_));
 sky130_vsdinv _32436_ (.A(_09727_),
    .Y(_10091_));
 sky130_fd_sc_hd__a21oi_4 _32437_ (.A1(_10089_),
    .A2(_10090_),
    .B1(_10091_),
    .Y(_10092_));
 sky130_vsdinv _32438_ (.A(_10079_),
    .Y(_10093_));
 sky130_fd_sc_hd__nand2_2 _32439_ (.A(_10088_),
    .B(_10076_),
    .Y(_10094_));
 sky130_fd_sc_hd__o211a_2 _32440_ (.A1(_10093_),
    .A2(_10094_),
    .B1(_10091_),
    .C1(_10089_),
    .X(_10095_));
 sky130_fd_sc_hd__o22ai_4 _32441_ (.A1(_10063_),
    .A2(_10064_),
    .B1(_10092_),
    .B2(_10095_),
    .Y(_10096_));
 sky130_fd_sc_hd__a21o_1 _32442_ (.A1(_10089_),
    .A2(_10090_),
    .B1(_10091_),
    .X(_10097_));
 sky130_fd_sc_hd__nand3_4 _32443_ (.A(_10089_),
    .B(_10091_),
    .C(_10090_),
    .Y(_10098_));
 sky130_fd_sc_hd__nand2_1 _32444_ (.A(_09687_),
    .B(_09700_),
    .Y(_10099_));
 sky130_fd_sc_hd__nand2_2 _32445_ (.A(_10099_),
    .B(_09683_),
    .Y(_10100_));
 sky130_fd_sc_hd__nand3_4 _32446_ (.A(_10097_),
    .B(_10098_),
    .C(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__nand2_2 _32447_ (.A(_10096_),
    .B(_10101_),
    .Y(_10102_));
 sky130_fd_sc_hd__nand2_2 _32448_ (.A(_10062_),
    .B(_10102_),
    .Y(_10103_));
 sky130_vsdinv _32449_ (.A(_09742_),
    .Y(_10104_));
 sky130_fd_sc_hd__nand2_1 _32450_ (.A(_09741_),
    .B(_10104_),
    .Y(_10105_));
 sky130_fd_sc_hd__nand2_1 _32451_ (.A(_10058_),
    .B(_10059_),
    .Y(_10106_));
 sky130_fd_sc_hd__o2111ai_4 _32452_ (.A1(_10054_),
    .A2(_10106_),
    .B1(_10096_),
    .C1(_10055_),
    .D1(_10101_),
    .Y(_10107_));
 sky130_fd_sc_hd__nand3_4 _32453_ (.A(_10103_),
    .B(_10105_),
    .C(_10107_),
    .Y(_10108_));
 sky130_fd_sc_hd__nand3_4 _32454_ (.A(_10062_),
    .B(_10096_),
    .C(_10101_),
    .Y(_10109_));
 sky130_fd_sc_hd__nand3_4 _32455_ (.A(_10102_),
    .B(_10055_),
    .C(_10061_),
    .Y(_10110_));
 sky130_fd_sc_hd__a31oi_4 _32456_ (.A1(_09707_),
    .A2(_09737_),
    .A3(_09740_),
    .B1(_09742_),
    .Y(_10111_));
 sky130_fd_sc_hd__nand3_4 _32457_ (.A(_10109_),
    .B(_10110_),
    .C(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__nand2_4 _32458_ (.A(_09643_),
    .B(_09645_),
    .Y(_10113_));
 sky130_fd_sc_hd__nand3_4 _32459_ (.A(_07743_),
    .B(_19634_),
    .C(_19893_),
    .Y(_10114_));
 sky130_fd_sc_hd__nor2_4 _32460_ (.A(_07274_),
    .B(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__nand2_2 _32461_ (.A(_06992_),
    .B(_06808_),
    .Y(_10116_));
 sky130_fd_sc_hd__a22o_1 _32462_ (.A1(_08190_),
    .A2(_06288_),
    .B1(_07928_),
    .B2(_06465_),
    .X(_10117_));
 sky130_fd_sc_hd__nand3b_2 _32463_ (.A_N(_10115_),
    .B(_10116_),
    .C(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__a21oi_4 _32464_ (.A1(_09690_),
    .A2(_09692_),
    .B1(_09697_),
    .Y(_10119_));
 sky130_fd_sc_hd__a22oi_4 _32465_ (.A1(_07744_),
    .A2(_06652_),
    .B1(_06921_),
    .B2(_07072_),
    .Y(_10120_));
 sky130_vsdinv _32466_ (.A(_10116_),
    .Y(_10121_));
 sky130_fd_sc_hd__o21ai_2 _32467_ (.A1(_10120_),
    .A2(_10115_),
    .B1(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__nand3_4 _32468_ (.A(_10118_),
    .B(_10119_),
    .C(_10122_),
    .Y(_10123_));
 sky130_fd_sc_hd__o21ai_2 _32469_ (.A1(_10120_),
    .A2(_10115_),
    .B1(_10116_),
    .Y(_10124_));
 sky130_fd_sc_hd__o21ai_2 _32470_ (.A1(_09691_),
    .A2(_09696_),
    .B1(_09689_),
    .Y(_10125_));
 sky130_fd_sc_hd__o211ai_4 _32471_ (.A1(net440),
    .A2(_10114_),
    .B1(_10121_),
    .C1(_10117_),
    .Y(_10126_));
 sky130_fd_sc_hd__nand3_4 _32472_ (.A(_10124_),
    .B(_10125_),
    .C(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__o21ai_4 _32473_ (.A1(_09631_),
    .A2(_09629_),
    .B1(_09636_),
    .Y(_10128_));
 sky130_fd_sc_hd__a21o_2 _32474_ (.A1(_10123_),
    .A2(_10127_),
    .B1(_10128_),
    .X(_10129_));
 sky130_fd_sc_hd__nand3_4 _32475_ (.A(_10123_),
    .B(_10127_),
    .C(_10128_),
    .Y(_10130_));
 sky130_fd_sc_hd__a22oi_4 _32476_ (.A1(_09639_),
    .A2(_10113_),
    .B1(_10129_),
    .B2(_10130_),
    .Y(_10131_));
 sky130_fd_sc_hd__nand2_1 _32477_ (.A(_09633_),
    .B(_09638_),
    .Y(_10132_));
 sky130_fd_sc_hd__o2111a_4 _32478_ (.A1(_09642_),
    .A2(_10132_),
    .B1(_10113_),
    .C1(_10130_),
    .D1(_10129_),
    .X(_10133_));
 sky130_fd_sc_hd__a22oi_4 _32479_ (.A1(_06341_),
    .A2(_07059_),
    .B1(_19647_),
    .B2(_08280_),
    .Y(_10134_));
 sky130_fd_sc_hd__nand2_4 _32480_ (.A(_19643_),
    .B(_19883_),
    .Y(_10135_));
 sky130_fd_sc_hd__nand2_4 _32481_ (.A(_19646_),
    .B(_06798_),
    .Y(_10136_));
 sky130_fd_sc_hd__nor2_4 _32482_ (.A(_10135_),
    .B(_10136_),
    .Y(_10137_));
 sky130_fd_sc_hd__nand2_2 _32483_ (.A(_06419_),
    .B(_19877_),
    .Y(_10138_));
 sky130_vsdinv _32484_ (.A(_10138_),
    .Y(_10139_));
 sky130_fd_sc_hd__o21ai_4 _32485_ (.A1(_10134_),
    .A2(_10137_),
    .B1(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__or2_1 _32486_ (.A(_10135_),
    .B(_10136_),
    .X(_10141_));
 sky130_fd_sc_hd__nand2_4 _32487_ (.A(_10135_),
    .B(_10136_),
    .Y(_10142_));
 sky130_fd_sc_hd__nand3_4 _32488_ (.A(_10141_),
    .B(_10138_),
    .C(_10142_),
    .Y(_10143_));
 sky130_fd_sc_hd__nor2_2 _32489_ (.A(_09616_),
    .B(_09614_),
    .Y(_10144_));
 sky130_fd_sc_hd__o2bb2ai_4 _32490_ (.A1_N(_10140_),
    .A2_N(_10143_),
    .B1(_09615_),
    .B2(_10144_),
    .Y(_10145_));
 sky130_fd_sc_hd__a21oi_2 _32491_ (.A1(_09619_),
    .A2(_09618_),
    .B1(_09615_),
    .Y(_10146_));
 sky130_fd_sc_hd__nand3_4 _32492_ (.A(_10143_),
    .B(_10146_),
    .C(_10140_),
    .Y(_10147_));
 sky130_fd_sc_hd__nand2_1 _32493_ (.A(_10145_),
    .B(_10147_),
    .Y(_10148_));
 sky130_fd_sc_hd__buf_4 _32494_ (.A(_08485_),
    .X(_10149_));
 sky130_fd_sc_hd__a22oi_4 _32495_ (.A1(_06326_),
    .A2(_19873_),
    .B1(_19654_),
    .B2(_07702_),
    .Y(_10150_));
 sky130_fd_sc_hd__nand2_2 _32496_ (.A(_06882_),
    .B(\pcpi_mul.rs1[18] ),
    .Y(_10151_));
 sky130_fd_sc_hd__nand2_2 _32497_ (.A(_05735_),
    .B(_07556_),
    .Y(_10152_));
 sky130_fd_sc_hd__nor2_4 _32498_ (.A(_10151_),
    .B(_10152_),
    .Y(_10153_));
 sky130_fd_sc_hd__a211o_1 _32499_ (.A1(_06014_),
    .A2(_10149_),
    .B1(_10150_),
    .C1(_10153_),
    .X(_10154_));
 sky130_fd_sc_hd__nand2_1 _32500_ (.A(_05731_),
    .B(_08485_),
    .Y(_10155_));
 sky130_vsdinv _32501_ (.A(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__o21ai_1 _32502_ (.A1(_10150_),
    .A2(_10153_),
    .B1(_10156_),
    .Y(_10157_));
 sky130_fd_sc_hd__nand2_2 _32503_ (.A(_10154_),
    .B(_10157_),
    .Y(_10158_));
 sky130_fd_sc_hd__nand2_1 _32504_ (.A(_10148_),
    .B(_10158_),
    .Y(_10159_));
 sky130_vsdinv _32505_ (.A(_10158_),
    .Y(_10160_));
 sky130_fd_sc_hd__nand3_1 _32506_ (.A(_10160_),
    .B(_10145_),
    .C(_10147_),
    .Y(_10161_));
 sky130_fd_sc_hd__nand2_2 _32507_ (.A(_10159_),
    .B(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__o21ai_2 _32508_ (.A1(_10131_),
    .A2(_10133_),
    .B1(_10162_),
    .Y(_10163_));
 sky130_fd_sc_hd__a21oi_2 _32509_ (.A1(_09738_),
    .A2(_09705_),
    .B1(_09704_),
    .Y(_10164_));
 sky130_fd_sc_hd__a22o_4 _32510_ (.A1(_09639_),
    .A2(_10113_),
    .B1(_10129_),
    .B2(_10130_),
    .X(_10165_));
 sky130_fd_sc_hd__nand2_1 _32511_ (.A(_10113_),
    .B(_09639_),
    .Y(_10166_));
 sky130_fd_sc_hd__nand3b_4 _32512_ (.A_N(_10166_),
    .B(_10130_),
    .C(_10129_),
    .Y(_10167_));
 sky130_fd_sc_hd__nand2_1 _32513_ (.A(_10148_),
    .B(_10160_),
    .Y(_10168_));
 sky130_fd_sc_hd__nand3_2 _32514_ (.A(_10145_),
    .B(_10158_),
    .C(_10147_),
    .Y(_10169_));
 sky130_fd_sc_hd__nand2_2 _32515_ (.A(_10168_),
    .B(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__nand3_2 _32516_ (.A(_10165_),
    .B(_10167_),
    .C(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__nand3_4 _32517_ (.A(_10163_),
    .B(_10164_),
    .C(_10171_),
    .Y(_10172_));
 sky130_vsdinv _32518_ (.A(_10169_),
    .Y(_10173_));
 sky130_fd_sc_hd__and2_1 _32519_ (.A(_10148_),
    .B(_10160_),
    .X(_10174_));
 sky130_fd_sc_hd__o22ai_4 _32520_ (.A1(_10173_),
    .A2(_10174_),
    .B1(_10131_),
    .B2(_10133_),
    .Y(_10175_));
 sky130_fd_sc_hd__o21ai_2 _32521_ (.A1(_09706_),
    .A2(_09703_),
    .B1(_09739_),
    .Y(_10176_));
 sky130_fd_sc_hd__nand3_4 _32522_ (.A(_10165_),
    .B(_10167_),
    .C(_10162_),
    .Y(_10177_));
 sky130_fd_sc_hd__nand3_4 _32523_ (.A(_10175_),
    .B(_10176_),
    .C(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__nand2_4 _32524_ (.A(_09659_),
    .B(_09655_),
    .Y(_10179_));
 sky130_fd_sc_hd__a21oi_1 _32525_ (.A1(_10172_),
    .A2(_10178_),
    .B1(_10179_),
    .Y(_10180_));
 sky130_fd_sc_hd__nand3_4 _32526_ (.A(_10172_),
    .B(_10178_),
    .C(_10179_),
    .Y(_10181_));
 sky130_vsdinv _32527_ (.A(_10181_),
    .Y(_10182_));
 sky130_fd_sc_hd__o2bb2ai_2 _32528_ (.A1_N(_10108_),
    .A2_N(_10112_),
    .B1(_10180_),
    .B2(_10182_),
    .Y(_10183_));
 sky130_fd_sc_hd__and3_2 _32529_ (.A(_10175_),
    .B(_10176_),
    .C(_10177_),
    .X(_10184_));
 sky130_fd_sc_hd__nand2_2 _32530_ (.A(_10172_),
    .B(_10179_),
    .Y(_10185_));
 sky130_fd_sc_hd__nand2_2 _32531_ (.A(_10172_),
    .B(_10178_),
    .Y(_10186_));
 sky130_vsdinv _32532_ (.A(_10179_),
    .Y(_10187_));
 sky130_fd_sc_hd__nand2_4 _32533_ (.A(_10186_),
    .B(_10187_),
    .Y(_10188_));
 sky130_fd_sc_hd__o2111ai_4 _32534_ (.A1(_10184_),
    .A2(_10185_),
    .B1(_10188_),
    .C1(_10108_),
    .D1(_10112_),
    .Y(_10189_));
 sky130_fd_sc_hd__nand3_4 _32535_ (.A(_10025_),
    .B(_10183_),
    .C(_10189_),
    .Y(_10190_));
 sky130_fd_sc_hd__nand2_1 _32536_ (.A(_10188_),
    .B(_10181_),
    .Y(_10191_));
 sky130_fd_sc_hd__nand3_4 _32537_ (.A(_10191_),
    .B(_10108_),
    .C(_10112_),
    .Y(_10192_));
 sky130_fd_sc_hd__a21oi_1 _32538_ (.A1(_10172_),
    .A2(_10178_),
    .B1(_10187_),
    .Y(_10193_));
 sky130_fd_sc_hd__nor2_1 _32539_ (.A(_10179_),
    .B(_10186_),
    .Y(_10194_));
 sky130_fd_sc_hd__o2bb2ai_2 _32540_ (.A1_N(_10108_),
    .A2_N(_10112_),
    .B1(_10193_),
    .B2(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__nor2_2 _32541_ (.A(_09751_),
    .B(_09754_),
    .Y(_10196_));
 sky130_fd_sc_hd__a31oi_4 _32542_ (.A1(_09663_),
    .A2(_09746_),
    .A3(_09671_),
    .B1(_10196_),
    .Y(_10197_));
 sky130_fd_sc_hd__nand3_4 _32543_ (.A(_10192_),
    .B(_10195_),
    .C(_10197_),
    .Y(_10198_));
 sky130_fd_sc_hd__nand3_4 _32544_ (.A(_10023_),
    .B(_10190_),
    .C(_10198_),
    .Y(_10199_));
 sky130_fd_sc_hd__a31oi_4 _32545_ (.A1(_09878_),
    .A2(_09872_),
    .A3(_09873_),
    .B1(_09762_),
    .Y(_10200_));
 sky130_fd_sc_hd__nand2_2 _32546_ (.A(_10198_),
    .B(_10190_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand3_4 _32547_ (.A(_10201_),
    .B(_10022_),
    .C(_10018_),
    .Y(_10202_));
 sky130_fd_sc_hd__nand3_4 _32548_ (.A(_10199_),
    .B(_10200_),
    .C(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__nand2_1 _32549_ (.A(_09758_),
    .B(_09755_),
    .Y(_10204_));
 sky130_fd_sc_hd__o22ai_4 _32550_ (.A1(_09875_),
    .A2(_10204_),
    .B1(_09759_),
    .B2(_09874_),
    .Y(_10205_));
 sky130_fd_sc_hd__a21oi_1 _32551_ (.A1(_10020_),
    .A2(_10021_),
    .B1(_10016_),
    .Y(_10206_));
 sky130_fd_sc_hd__nor3_4 _32552_ (.A(_10017_),
    .B(_10012_),
    .C(_10014_),
    .Y(_10207_));
 sky130_fd_sc_hd__o21ai_2 _32553_ (.A1(_10206_),
    .A2(_10207_),
    .B1(_10201_),
    .Y(_10208_));
 sky130_fd_sc_hd__nand2_2 _32554_ (.A(_10020_),
    .B(_10016_),
    .Y(_10209_));
 sky130_fd_sc_hd__o2111ai_4 _32555_ (.A1(_10014_),
    .A2(_10209_),
    .B1(_10190_),
    .C1(_10198_),
    .D1(_10018_),
    .Y(_10210_));
 sky130_fd_sc_hd__nand3_4 _32556_ (.A(_10205_),
    .B(_10208_),
    .C(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__nand2_1 _32557_ (.A(_10203_),
    .B(_10211_),
    .Y(_10212_));
 sky130_fd_sc_hd__nor2_4 _32558_ (.A(_09871_),
    .B(_09857_),
    .Y(_10213_));
 sky130_vsdinv _32559_ (.A(_09840_),
    .Y(_10214_));
 sky130_fd_sc_hd__a21oi_4 _32560_ (.A1(_09843_),
    .A2(_09836_),
    .B1(_10214_),
    .Y(_10215_));
 sky130_fd_sc_hd__nand2_1 _32561_ (.A(_10213_),
    .B(_10215_),
    .Y(_10216_));
 sky130_fd_sc_hd__a21o_1 _32562_ (.A1(_09884_),
    .A2(_09853_),
    .B1(_10215_),
    .X(_10217_));
 sky130_fd_sc_hd__nand2_2 _32563_ (.A(_10216_),
    .B(_10217_),
    .Y(_10218_));
 sky130_vsdinv _32564_ (.A(_10218_),
    .Y(_10219_));
 sky130_fd_sc_hd__nand2_1 _32565_ (.A(_10212_),
    .B(_10219_),
    .Y(_10220_));
 sky130_fd_sc_hd__nand3_2 _32566_ (.A(_10203_),
    .B(_10211_),
    .C(_10218_),
    .Y(_10221_));
 sky130_fd_sc_hd__a21boi_4 _32567_ (.A1(_09881_),
    .A2(_09897_),
    .B1_N(_09888_),
    .Y(_10222_));
 sky130_fd_sc_hd__nand3_2 _32568_ (.A(_10220_),
    .B(_10221_),
    .C(_10222_),
    .Y(_10223_));
 sky130_vsdinv _32569_ (.A(_10217_),
    .Y(_10224_));
 sky130_fd_sc_hd__and3_1 _32570_ (.A(_09884_),
    .B(_09853_),
    .C(_10215_),
    .X(_10225_));
 sky130_fd_sc_hd__o2bb2ai_2 _32571_ (.A1_N(_10211_),
    .A2_N(_10203_),
    .B1(_10224_),
    .B2(_10225_),
    .Y(_10226_));
 sky130_vsdinv _32572_ (.A(_09883_),
    .Y(_10227_));
 sky130_fd_sc_hd__nand2_1 _32573_ (.A(_09887_),
    .B(_09885_),
    .Y(_10228_));
 sky130_fd_sc_hd__o2bb2ai_2 _32574_ (.A1_N(_09881_),
    .A2_N(_09897_),
    .B1(_10227_),
    .B2(_10228_),
    .Y(_10229_));
 sky130_fd_sc_hd__nand3_2 _32575_ (.A(_10219_),
    .B(_10203_),
    .C(_10211_),
    .Y(_10230_));
 sky130_fd_sc_hd__nand3_4 _32576_ (.A(_10226_),
    .B(_10229_),
    .C(_10230_),
    .Y(_10231_));
 sky130_fd_sc_hd__nand2_1 _32577_ (.A(_10223_),
    .B(_10231_),
    .Y(_10232_));
 sky130_vsdinv _32578_ (.A(_09896_),
    .Y(_10233_));
 sky130_fd_sc_hd__nand2_1 _32579_ (.A(_10232_),
    .B(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__a31oi_2 _32580_ (.A1(_10220_),
    .A2(_10222_),
    .A3(_10221_),
    .B1(_10233_),
    .Y(_10235_));
 sky130_fd_sc_hd__nand2_1 _32581_ (.A(_10235_),
    .B(_10231_),
    .Y(_10236_));
 sky130_fd_sc_hd__nand3b_4 _32582_ (.A_N(_09926_),
    .B(_10234_),
    .C(_10236_),
    .Y(_10237_));
 sky130_fd_sc_hd__nand2_1 _32583_ (.A(_10232_),
    .B(_09896_),
    .Y(_10238_));
 sky130_fd_sc_hd__nand3_2 _32584_ (.A(_10223_),
    .B(_10231_),
    .C(_10233_),
    .Y(_10239_));
 sky130_fd_sc_hd__nand3_4 _32585_ (.A(_10238_),
    .B(_10239_),
    .C(_09926_),
    .Y(_10240_));
 sky130_fd_sc_hd__nand2_2 _32586_ (.A(_10237_),
    .B(_10240_),
    .Y(_10241_));
 sky130_fd_sc_hd__nand2_1 _32587_ (.A(_09925_),
    .B(_09915_),
    .Y(_10242_));
 sky130_fd_sc_hd__nand2_2 _32588_ (.A(_10242_),
    .B(_09917_),
    .Y(_10243_));
 sky130_fd_sc_hd__xor2_4 _32589_ (.A(_10241_),
    .B(_10243_),
    .X(_02648_));
 sky130_fd_sc_hd__a21oi_4 _32590_ (.A1(_10199_),
    .A2(_10202_),
    .B1(_10200_),
    .Y(_10244_));
 sky130_fd_sc_hd__a31oi_4 _32591_ (.A1(_10199_),
    .A2(_10200_),
    .A3(_10202_),
    .B1(_10218_),
    .Y(_10245_));
 sky130_fd_sc_hd__nand3_1 _32592_ (.A(_10018_),
    .B(_10022_),
    .C(_10198_),
    .Y(_10246_));
 sky130_fd_sc_hd__nand2_2 _32593_ (.A(_10246_),
    .B(_10190_),
    .Y(_10247_));
 sky130_fd_sc_hd__a21oi_4 _32594_ (.A1(_10109_),
    .A2(_10110_),
    .B1(_10111_),
    .Y(_10248_));
 sky130_fd_sc_hd__a31oi_4 _32595_ (.A1(_10112_),
    .A2(_10188_),
    .A3(_10181_),
    .B1(_10248_),
    .Y(_10249_));
 sky130_fd_sc_hd__nand2_2 _32596_ (.A(_10047_),
    .B(_10048_),
    .Y(_10250_));
 sky130_fd_sc_hd__buf_6 _32597_ (.A(\pcpi_mul.rs2[27] ),
    .X(_10251_));
 sky130_fd_sc_hd__a31o_1 _32598_ (.A1(_10250_),
    .A2(_10251_),
    .A3(_19928_),
    .B1(_10049_),
    .X(_10252_));
 sky130_fd_sc_hd__nor2_4 _32599_ (.A(_09509_),
    .B(_10026_),
    .Y(_10253_));
 sky130_fd_sc_hd__nand2_2 _32600_ (.A(_19602_),
    .B(_19913_),
    .Y(_10254_));
 sky130_vsdinv _32601_ (.A(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__clkbuf_4 _32602_ (.A(\pcpi_mul.rs2[26] ),
    .X(_10256_));
 sky130_fd_sc_hd__buf_4 _32603_ (.A(_08945_),
    .X(_10257_));
 sky130_fd_sc_hd__a22o_2 _32604_ (.A1(_10256_),
    .A2(_05374_),
    .B1(_10257_),
    .B2(_19917_),
    .X(_10258_));
 sky130_fd_sc_hd__nand3b_4 _32605_ (.A_N(_10253_),
    .B(_10255_),
    .C(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__buf_6 _32606_ (.A(_19595_),
    .X(_10260_));
 sky130_fd_sc_hd__buf_4 _32607_ (.A(_19599_),
    .X(_10261_));
 sky130_fd_sc_hd__a22oi_4 _32608_ (.A1(_10260_),
    .A2(_05174_),
    .B1(_10261_),
    .B2(_05493_),
    .Y(_10262_));
 sky130_fd_sc_hd__o21ai_2 _32609_ (.A1(_10262_),
    .A2(_10253_),
    .B1(_10254_),
    .Y(_10263_));
 sky130_fd_sc_hd__nand3_4 _32610_ (.A(_10252_),
    .B(_10259_),
    .C(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__a21oi_4 _32611_ (.A1(_10045_),
    .A2(_10250_),
    .B1(_10049_),
    .Y(_10265_));
 sky130_fd_sc_hd__o21ai_2 _32612_ (.A1(_10262_),
    .A2(_10253_),
    .B1(_10255_),
    .Y(_10266_));
 sky130_fd_sc_hd__o211ai_4 _32613_ (.A1(_09509_),
    .A2(_10026_),
    .B1(_10254_),
    .C1(_10258_),
    .Y(_10267_));
 sky130_fd_sc_hd__nand3_2 _32614_ (.A(_10265_),
    .B(_10266_),
    .C(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__o21ai_2 _32615_ (.A1(_10033_),
    .A2(_10027_),
    .B1(_10029_),
    .Y(_10269_));
 sky130_vsdinv _32616_ (.A(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__a21o_2 _32617_ (.A1(_10264_),
    .A2(_10268_),
    .B1(_10270_),
    .X(_10271_));
 sky130_fd_sc_hd__a31oi_4 _32618_ (.A1(_10265_),
    .A2(_10266_),
    .A3(_10267_),
    .B1(_10269_),
    .Y(_10272_));
 sky130_fd_sc_hd__nand2_2 _32619_ (.A(_10272_),
    .B(_10264_),
    .Y(_10273_));
 sky130_fd_sc_hd__nand2_2 _32620_ (.A(_19582_),
    .B(_05122_),
    .Y(_10274_));
 sky130_fd_sc_hd__nand2_2 _32621_ (.A(_19586_),
    .B(_07828_),
    .Y(_10275_));
 sky130_fd_sc_hd__or2_1 _32622_ (.A(_10274_),
    .B(_10275_),
    .X(_10276_));
 sky130_fd_sc_hd__nand2_2 _32623_ (.A(_10274_),
    .B(_10275_),
    .Y(_10277_));
 sky130_fd_sc_hd__nand2_2 _32624_ (.A(_19591_),
    .B(_05467_),
    .Y(_10278_));
 sky130_vsdinv _32625_ (.A(_10278_),
    .Y(_10279_));
 sky130_fd_sc_hd__nand3_4 _32626_ (.A(_10276_),
    .B(_10277_),
    .C(_10279_),
    .Y(_10280_));
 sky130_fd_sc_hd__buf_4 _32627_ (.A(_19582_),
    .X(_10281_));
 sky130_fd_sc_hd__buf_6 _32628_ (.A(_19586_),
    .X(_10282_));
 sky130_fd_sc_hd__a22oi_4 _32629_ (.A1(_10281_),
    .A2(_07759_),
    .B1(_10282_),
    .B2(_05230_),
    .Y(_10283_));
 sky130_fd_sc_hd__nor2_2 _32630_ (.A(_10274_),
    .B(_10275_),
    .Y(_10284_));
 sky130_fd_sc_hd__o21ai_2 _32631_ (.A1(_10283_),
    .A2(_10284_),
    .B1(_10278_),
    .Y(_10285_));
 sky130_fd_sc_hd__clkinv_8 _32632_ (.A(net498),
    .Y(_10286_));
 sky130_fd_sc_hd__nor2_4 _32633_ (.A(_10286_),
    .B(_04841_),
    .Y(_10287_));
 sky130_fd_sc_hd__a21o_1 _32634_ (.A1(_10280_),
    .A2(_10285_),
    .B1(_10287_),
    .X(_10288_));
 sky130_fd_sc_hd__nand3_4 _32635_ (.A(_10280_),
    .B(_10287_),
    .C(_10285_),
    .Y(_10289_));
 sky130_fd_sc_hd__nand2_2 _32636_ (.A(_10288_),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__a21boi_4 _32637_ (.A1(_10271_),
    .A2(_10273_),
    .B1_N(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__nand2_1 _32638_ (.A(_10268_),
    .B(_10270_),
    .Y(_10292_));
 sky130_fd_sc_hd__and3_2 _32639_ (.A(_10252_),
    .B(_10259_),
    .C(_10263_),
    .X(_10293_));
 sky130_fd_sc_hd__o2111a_4 _32640_ (.A1(_10292_),
    .A2(_10293_),
    .B1(_10288_),
    .C1(_10289_),
    .D1(_10271_),
    .X(_10294_));
 sky130_fd_sc_hd__o22ai_4 _32641_ (.A1(_10057_),
    .A2(_10056_),
    .B1(_10291_),
    .B2(_10294_),
    .Y(_10295_));
 sky130_fd_sc_hd__nand2_2 _32642_ (.A(_10271_),
    .B(_10273_),
    .Y(_10296_));
 sky130_fd_sc_hd__nand2_1 _32643_ (.A(_10296_),
    .B(_10290_),
    .Y(_10297_));
 sky130_fd_sc_hd__nand3b_2 _32644_ (.A_N(_10290_),
    .B(_10271_),
    .C(_10273_),
    .Y(_10298_));
 sky130_fd_sc_hd__nand3_4 _32645_ (.A(_10297_),
    .B(_10054_),
    .C(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__nand2_2 _32646_ (.A(_10295_),
    .B(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__nand3_4 _32647_ (.A(_09191_),
    .B(_19610_),
    .C(_19909_),
    .Y(_10301_));
 sky130_fd_sc_hd__nor2_8 _32648_ (.A(_05663_),
    .B(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__nand2_4 _32649_ (.A(_08545_),
    .B(_06826_),
    .Y(_10303_));
 sky130_vsdinv _32650_ (.A(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__a22o_2 _32651_ (.A1(_08549_),
    .A2(_08198_),
    .B1(_09680_),
    .B2(_05661_),
    .X(_10305_));
 sky130_fd_sc_hd__nand3b_2 _32652_ (.A_N(_10302_),
    .B(_10304_),
    .C(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__o22ai_4 _32653_ (.A1(_06215_),
    .A2(_10068_),
    .B1(_10070_),
    .B2(_10067_),
    .Y(_10307_));
 sky130_fd_sc_hd__a22oi_4 _32654_ (.A1(_08152_),
    .A2(_05545_),
    .B1(_07984_),
    .B2(_06105_),
    .Y(_10308_));
 sky130_fd_sc_hd__o21ai_2 _32655_ (.A1(_10308_),
    .A2(_10302_),
    .B1(_10303_),
    .Y(_10309_));
 sky130_fd_sc_hd__nand3_4 _32656_ (.A(_10306_),
    .B(_10307_),
    .C(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__o21ai_2 _32657_ (.A1(_10308_),
    .A2(_10302_),
    .B1(_10304_),
    .Y(_10311_));
 sky130_fd_sc_hd__a21oi_2 _32658_ (.A1(_10074_),
    .A2(_10071_),
    .B1(_10069_),
    .Y(_10312_));
 sky130_fd_sc_hd__o211ai_4 _32659_ (.A1(_08189_),
    .A2(_10301_),
    .B1(_10303_),
    .C1(_10305_),
    .Y(_10313_));
 sky130_fd_sc_hd__nand3_4 _32660_ (.A(_10311_),
    .B(_10312_),
    .C(_10313_),
    .Y(_10314_));
 sky130_fd_sc_hd__nand2_1 _32661_ (.A(_10310_),
    .B(_10314_),
    .Y(_10315_));
 sky130_fd_sc_hd__nand2_2 _32662_ (.A(_07933_),
    .B(_06259_),
    .Y(_10316_));
 sky130_fd_sc_hd__nand2_2 _32663_ (.A(_07824_),
    .B(_06648_),
    .Y(_10317_));
 sky130_fd_sc_hd__nor2_4 _32664_ (.A(_10316_),
    .B(_10317_),
    .Y(_10318_));
 sky130_fd_sc_hd__and2_1 _32665_ (.A(_10316_),
    .B(_10317_),
    .X(_10319_));
 sky130_fd_sc_hd__nand2_2 _32666_ (.A(_19627_),
    .B(_19894_),
    .Y(_10320_));
 sky130_vsdinv _32667_ (.A(_10320_),
    .Y(_10321_));
 sky130_fd_sc_hd__o21ai_4 _32668_ (.A1(_10318_),
    .A2(_10319_),
    .B1(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__nand2_2 _32669_ (.A(_10316_),
    .B(_10317_),
    .Y(_10323_));
 sky130_fd_sc_hd__nand3b_4 _32670_ (.A_N(_10318_),
    .B(_10323_),
    .C(_10320_),
    .Y(_10324_));
 sky130_fd_sc_hd__and2_1 _32671_ (.A(_10322_),
    .B(_10324_),
    .X(_10325_));
 sky130_fd_sc_hd__nand2_4 _32672_ (.A(_10315_),
    .B(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__nand2_2 _32673_ (.A(_10322_),
    .B(_10324_),
    .Y(_10327_));
 sky130_fd_sc_hd__nand3_4 _32674_ (.A(_10327_),
    .B(_10310_),
    .C(_10314_),
    .Y(_10328_));
 sky130_vsdinv _32675_ (.A(_10040_),
    .Y(_10329_));
 sky130_fd_sc_hd__nand2_1 _32676_ (.A(_10035_),
    .B(_10329_),
    .Y(_10330_));
 sky130_fd_sc_hd__nand2_2 _32677_ (.A(_10330_),
    .B(_10038_),
    .Y(_10331_));
 sky130_fd_sc_hd__a21oi_2 _32678_ (.A1(_10326_),
    .A2(_10328_),
    .B1(_10331_),
    .Y(_10332_));
 sky130_vsdinv _32679_ (.A(_10038_),
    .Y(_10333_));
 sky130_fd_sc_hd__o211a_4 _32680_ (.A1(_10042_),
    .A2(_10333_),
    .B1(_10328_),
    .C1(_10326_),
    .X(_10334_));
 sky130_fd_sc_hd__nand2_4 _32681_ (.A(_10094_),
    .B(_10079_),
    .Y(_10335_));
 sky130_fd_sc_hd__o21bai_4 _32682_ (.A1(_10332_),
    .A2(_10334_),
    .B1_N(_10335_),
    .Y(_10336_));
 sky130_vsdinv _32683_ (.A(_10035_),
    .Y(_10337_));
 sky130_fd_sc_hd__and2_1 _32684_ (.A(_10038_),
    .B(_10040_),
    .X(_10338_));
 sky130_fd_sc_hd__o2bb2ai_4 _32685_ (.A1_N(_10328_),
    .A2_N(_10326_),
    .B1(_10337_),
    .B2(_10338_),
    .Y(_10339_));
 sky130_fd_sc_hd__nand3_4 _32686_ (.A(_10326_),
    .B(_10331_),
    .C(_10328_),
    .Y(_10340_));
 sky130_fd_sc_hd__nand3_4 _32687_ (.A(_10339_),
    .B(_10340_),
    .C(_10335_),
    .Y(_10341_));
 sky130_fd_sc_hd__nand3_4 _32688_ (.A(_10300_),
    .B(_10336_),
    .C(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__nor3_4 _32689_ (.A(_09734_),
    .B(_10053_),
    .C(_10054_),
    .Y(_10343_));
 sky130_fd_sc_hd__a31oi_4 _32690_ (.A1(_10055_),
    .A2(_10096_),
    .A3(_10101_),
    .B1(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__nand2_2 _32691_ (.A(_10336_),
    .B(_10341_),
    .Y(_10345_));
 sky130_fd_sc_hd__nand3_4 _32692_ (.A(_10345_),
    .B(_10295_),
    .C(_10299_),
    .Y(_10346_));
 sky130_fd_sc_hd__nand3_4 _32693_ (.A(_10342_),
    .B(_10344_),
    .C(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__a31o_1 _32694_ (.A1(_10055_),
    .A2(_10096_),
    .A3(_10101_),
    .B1(_10343_),
    .X(_10348_));
 sky130_fd_sc_hd__nand2_4 _32695_ (.A(_10300_),
    .B(_10345_),
    .Y(_10349_));
 sky130_fd_sc_hd__nand2_2 _32696_ (.A(_10339_),
    .B(_10335_),
    .Y(_10350_));
 sky130_fd_sc_hd__o2111ai_4 _32697_ (.A1(_10334_),
    .A2(_10350_),
    .B1(_10299_),
    .C1(_10336_),
    .D1(_10295_),
    .Y(_10351_));
 sky130_fd_sc_hd__nand3_4 _32698_ (.A(_10348_),
    .B(_10349_),
    .C(_10351_),
    .Y(_10352_));
 sky130_fd_sc_hd__nor2_2 _32699_ (.A(_10100_),
    .B(_10095_),
    .Y(_10353_));
 sky130_vsdinv _32700_ (.A(_10123_),
    .Y(_10354_));
 sky130_fd_sc_hd__a31o_1 _32701_ (.A1(_10124_),
    .A2(_10125_),
    .A3(_10126_),
    .B1(_10128_),
    .X(_10355_));
 sky130_vsdinv _32702_ (.A(_10355_),
    .Y(_10356_));
 sky130_fd_sc_hd__nand2_4 _32703_ (.A(_06923_),
    .B(_19890_),
    .Y(_10357_));
 sky130_fd_sc_hd__nand2_4 _32704_ (.A(_06920_),
    .B(_06808_),
    .Y(_10358_));
 sky130_fd_sc_hd__nor2_8 _32705_ (.A(_10357_),
    .B(_10358_),
    .Y(_10359_));
 sky130_fd_sc_hd__and2_2 _32706_ (.A(_10357_),
    .B(_10358_),
    .X(_10360_));
 sky130_fd_sc_hd__nand2_2 _32707_ (.A(_19641_),
    .B(_06443_),
    .Y(_10361_));
 sky130_fd_sc_hd__o21ai_2 _32708_ (.A1(_10359_),
    .A2(_10360_),
    .B1(_10361_),
    .Y(_10362_));
 sky130_fd_sc_hd__nand2_1 _32709_ (.A(_10081_),
    .B(_10082_),
    .Y(_10363_));
 sky130_fd_sc_hd__buf_4 _32710_ (.A(_07481_),
    .X(_10364_));
 sky130_fd_sc_hd__buf_4 _32711_ (.A(_06657_),
    .X(_10365_));
 sky130_fd_sc_hd__a31o_1 _32712_ (.A1(_10363_),
    .A2(_10364_),
    .A3(_10365_),
    .B1(_10083_),
    .X(_10366_));
 sky130_vsdinv _32713_ (.A(_10361_),
    .Y(_10367_));
 sky130_fd_sc_hd__nand2_2 _32714_ (.A(_10357_),
    .B(_10358_),
    .Y(_10368_));
 sky130_fd_sc_hd__nand3b_2 _32715_ (.A_N(_10359_),
    .B(_10367_),
    .C(_10368_),
    .Y(_10369_));
 sky130_fd_sc_hd__nand3_4 _32716_ (.A(_10362_),
    .B(_10366_),
    .C(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__o21ai_2 _32717_ (.A1(_10359_),
    .A2(_10360_),
    .B1(_10367_),
    .Y(_10371_));
 sky130_fd_sc_hd__nand3b_2 _32718_ (.A_N(_10359_),
    .B(_10361_),
    .C(_10368_),
    .Y(_10372_));
 sky130_fd_sc_hd__a21oi_2 _32719_ (.A1(_10086_),
    .A2(_10363_),
    .B1(_10083_),
    .Y(_10373_));
 sky130_fd_sc_hd__nand3_4 _32720_ (.A(_10371_),
    .B(_10372_),
    .C(_10373_),
    .Y(_10374_));
 sky130_fd_sc_hd__o21a_2 _32721_ (.A1(_10121_),
    .A2(_10115_),
    .B1(_10117_),
    .X(_10375_));
 sky130_fd_sc_hd__a21oi_4 _32722_ (.A1(_10370_),
    .A2(_10374_),
    .B1(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__and3_1 _32723_ (.A(_10370_),
    .B(_10374_),
    .C(_10375_),
    .X(_10377_));
 sky130_fd_sc_hd__o22ai_4 _32724_ (.A1(_10354_),
    .A2(_10356_),
    .B1(_10376_),
    .B2(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__a21o_1 _32725_ (.A1(_10370_),
    .A2(_10374_),
    .B1(_10375_),
    .X(_10379_));
 sky130_fd_sc_hd__nand2_2 _32726_ (.A(_10130_),
    .B(_10127_),
    .Y(_10380_));
 sky130_fd_sc_hd__nand3_4 _32727_ (.A(_10370_),
    .B(_10374_),
    .C(_10375_),
    .Y(_10381_));
 sky130_fd_sc_hd__nand3_4 _32728_ (.A(_10379_),
    .B(_10380_),
    .C(_10381_),
    .Y(_10382_));
 sky130_fd_sc_hd__nand2_4 _32729_ (.A(_06608_),
    .B(_06654_),
    .Y(_10383_));
 sky130_fd_sc_hd__nand2_4 _32730_ (.A(_06610_),
    .B(_19877_),
    .Y(_10384_));
 sky130_fd_sc_hd__nor2_8 _32731_ (.A(_10383_),
    .B(_10384_),
    .Y(_10385_));
 sky130_fd_sc_hd__and2_1 _32732_ (.A(_10383_),
    .B(_10384_),
    .X(_10386_));
 sky130_fd_sc_hd__nand2_2 _32733_ (.A(_06349_),
    .B(_07346_),
    .Y(_10387_));
 sky130_fd_sc_hd__o21bai_2 _32734_ (.A1(_10385_),
    .A2(_10386_),
    .B1_N(_10387_),
    .Y(_10388_));
 sky130_fd_sc_hd__nand2_2 _32735_ (.A(_10383_),
    .B(_10384_),
    .Y(_10389_));
 sky130_fd_sc_hd__nand3b_4 _32736_ (.A_N(_10385_),
    .B(_10387_),
    .C(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__a21oi_4 _32737_ (.A1(_10139_),
    .A2(_10142_),
    .B1(_10137_),
    .Y(_10391_));
 sky130_fd_sc_hd__nand3_4 _32738_ (.A(_10388_),
    .B(_10390_),
    .C(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__a21o_2 _32739_ (.A1(_10388_),
    .A2(_10390_),
    .B1(_10391_),
    .X(_10393_));
 sky130_fd_sc_hd__buf_6 _32740_ (.A(_07556_),
    .X(_10394_));
 sky130_fd_sc_hd__buf_6 _32741_ (.A(_07542_),
    .X(_10395_));
 sky130_fd_sc_hd__a22oi_4 _32742_ (.A1(_06883_),
    .A2(_10394_),
    .B1(_06884_),
    .B2(_10395_),
    .Y(_10396_));
 sky130_fd_sc_hd__nand3_4 _32743_ (.A(_06018_),
    .B(_06024_),
    .C(_07325_),
    .Y(_10397_));
 sky130_fd_sc_hd__nor2_1 _32744_ (.A(_08079_),
    .B(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__nand2_2 _32745_ (.A(_19659_),
    .B(_09772_),
    .Y(_10399_));
 sky130_fd_sc_hd__o21bai_1 _32746_ (.A1(_10396_),
    .A2(_10398_),
    .B1_N(_10399_),
    .Y(_10400_));
 sky130_vsdinv _32747_ (.A(_10400_),
    .Y(_10401_));
 sky130_fd_sc_hd__nor2_1 _32748_ (.A(_10396_),
    .B(_10398_),
    .Y(_10402_));
 sky130_fd_sc_hd__nand2_1 _32749_ (.A(_10402_),
    .B(_10399_),
    .Y(_10403_));
 sky130_vsdinv _32750_ (.A(_10403_),
    .Y(_10404_));
 sky130_fd_sc_hd__o2bb2ai_4 _32751_ (.A1_N(_10392_),
    .A2_N(_10393_),
    .B1(_10401_),
    .B2(_10404_),
    .Y(_10405_));
 sky130_fd_sc_hd__nand2_2 _32752_ (.A(_10403_),
    .B(_10400_),
    .Y(_10406_));
 sky130_fd_sc_hd__nand3b_4 _32753_ (.A_N(_10406_),
    .B(_10393_),
    .C(_10392_),
    .Y(_10407_));
 sky130_fd_sc_hd__nand2_8 _32754_ (.A(_10405_),
    .B(_10407_),
    .Y(_10408_));
 sky130_fd_sc_hd__a21oi_2 _32755_ (.A1(_10378_),
    .A2(_10382_),
    .B1(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__nand3_4 _32756_ (.A(_10381_),
    .B(_10123_),
    .C(_10355_),
    .Y(_10410_));
 sky130_fd_sc_hd__o211a_1 _32757_ (.A1(_10376_),
    .A2(_10410_),
    .B1(_10408_),
    .C1(_10378_),
    .X(_10411_));
 sky130_fd_sc_hd__o22ai_4 _32758_ (.A1(_10092_),
    .A2(_10353_),
    .B1(_10409_),
    .B2(_10411_),
    .Y(_10412_));
 sky130_fd_sc_hd__nor2_8 _32759_ (.A(_10376_),
    .B(_10410_),
    .Y(_10413_));
 sky130_fd_sc_hd__a21oi_4 _32760_ (.A1(_10379_),
    .A2(_10381_),
    .B1(_10380_),
    .Y(_10414_));
 sky130_fd_sc_hd__o21bai_4 _32761_ (.A1(_10413_),
    .A2(_10414_),
    .B1_N(_10408_),
    .Y(_10415_));
 sky130_vsdinv _32762_ (.A(_10100_),
    .Y(_10416_));
 sky130_fd_sc_hd__o21ai_4 _32763_ (.A1(_10416_),
    .A2(_10092_),
    .B1(_10098_),
    .Y(_10417_));
 sky130_fd_sc_hd__nand3_4 _32764_ (.A(_10378_),
    .B(_10408_),
    .C(_10382_),
    .Y(_10418_));
 sky130_fd_sc_hd__nand3_4 _32765_ (.A(_10415_),
    .B(_10417_),
    .C(_10418_),
    .Y(_10419_));
 sky130_fd_sc_hd__nand2_2 _32766_ (.A(_10170_),
    .B(_10167_),
    .Y(_10420_));
 sky130_fd_sc_hd__nand2_4 _32767_ (.A(_10420_),
    .B(_10165_),
    .Y(_10421_));
 sky130_fd_sc_hd__a21oi_2 _32768_ (.A1(_10412_),
    .A2(_10419_),
    .B1(_10421_),
    .Y(_10422_));
 sky130_fd_sc_hd__a21oi_4 _32769_ (.A1(_10415_),
    .A2(_10418_),
    .B1(_10417_),
    .Y(_10423_));
 sky130_fd_sc_hd__nand2_2 _32770_ (.A(_10419_),
    .B(_10421_),
    .Y(_10424_));
 sky130_fd_sc_hd__nor2_2 _32771_ (.A(_10423_),
    .B(_10424_),
    .Y(_10425_));
 sky130_fd_sc_hd__o2bb2ai_4 _32772_ (.A1_N(_10347_),
    .A2_N(_10352_),
    .B1(_10422_),
    .B2(_10425_),
    .Y(_10426_));
 sky130_fd_sc_hd__nor2_1 _32773_ (.A(_10416_),
    .B(_10092_),
    .Y(_10427_));
 sky130_fd_sc_hd__o211a_4 _32774_ (.A1(_10095_),
    .A2(_10427_),
    .B1(_10418_),
    .C1(_10415_),
    .X(_10428_));
 sky130_vsdinv _32775_ (.A(_10421_),
    .Y(_10429_));
 sky130_fd_sc_hd__o21ai_2 _32776_ (.A1(_10423_),
    .A2(_10428_),
    .B1(_10429_),
    .Y(_10430_));
 sky130_fd_sc_hd__o2111ai_4 _32777_ (.A1(_10423_),
    .A2(_10424_),
    .B1(_10347_),
    .C1(_10352_),
    .D1(_10430_),
    .Y(_10431_));
 sky130_fd_sc_hd__nand3_4 _32778_ (.A(_10249_),
    .B(_10426_),
    .C(_10431_),
    .Y(_10432_));
 sky130_fd_sc_hd__nand3_1 _32779_ (.A(_10112_),
    .B(_10188_),
    .C(_10181_),
    .Y(_10433_));
 sky130_fd_sc_hd__nand2_1 _32780_ (.A(_10433_),
    .B(_10108_),
    .Y(_10434_));
 sky130_fd_sc_hd__a21oi_1 _32781_ (.A1(_10412_),
    .A2(_10419_),
    .B1(_10429_),
    .Y(_10435_));
 sky130_fd_sc_hd__nor2_1 _32782_ (.A(_10131_),
    .B(_10170_),
    .Y(_10436_));
 sky130_fd_sc_hd__o211a_1 _32783_ (.A1(_10133_),
    .A2(_10436_),
    .B1(_10419_),
    .C1(_10412_),
    .X(_10437_));
 sky130_fd_sc_hd__o2bb2ai_2 _32784_ (.A1_N(_10347_),
    .A2_N(_10352_),
    .B1(_10435_),
    .B2(_10437_),
    .Y(_10438_));
 sky130_fd_sc_hd__nand2_1 _32785_ (.A(_10412_),
    .B(_10429_),
    .Y(_10439_));
 sky130_vsdinv _32786_ (.A(_10420_),
    .Y(_10440_));
 sky130_fd_sc_hd__o22ai_4 _32787_ (.A1(_10131_),
    .A2(_10440_),
    .B1(_10423_),
    .B2(_10428_),
    .Y(_10441_));
 sky130_fd_sc_hd__o2111ai_4 _32788_ (.A1(_10428_),
    .A2(_10439_),
    .B1(_10347_),
    .C1(_10352_),
    .D1(_10441_),
    .Y(_10442_));
 sky130_fd_sc_hd__nand3_4 _32789_ (.A(_10434_),
    .B(_10438_),
    .C(_10442_),
    .Y(_10443_));
 sky130_fd_sc_hd__nand2_1 _32790_ (.A(_10432_),
    .B(_10443_),
    .Y(_10444_));
 sky130_vsdinv _32791_ (.A(_09998_),
    .Y(_10445_));
 sky130_fd_sc_hd__nand2_1 _32792_ (.A(_09997_),
    .B(_10445_),
    .Y(_10446_));
 sky130_vsdinv _32793_ (.A(_09979_),
    .Y(_10447_));
 sky130_fd_sc_hd__nor2_2 _32794_ (.A(_09984_),
    .B(_09990_),
    .Y(_10448_));
 sky130_vsdinv _32795_ (.A(\pcpi_mul.rs1[23] ),
    .Y(_10449_));
 sky130_fd_sc_hd__nand3_4 _32796_ (.A(_05591_),
    .B(_19664_),
    .C(_08331_),
    .Y(_10450_));
 sky130_fd_sc_hd__nor2_4 _32797_ (.A(_10449_),
    .B(_10450_),
    .Y(_10451_));
 sky130_fd_sc_hd__nand2_2 _32798_ (.A(_19667_),
    .B(_09076_),
    .Y(_10452_));
 sky130_fd_sc_hd__clkbuf_4 _32799_ (.A(_09972_),
    .X(_10453_));
 sky130_fd_sc_hd__a22o_2 _32800_ (.A1(_06076_),
    .A2(_08337_),
    .B1(_06835_),
    .B2(_10453_),
    .X(_10454_));
 sky130_fd_sc_hd__nand3b_2 _32801_ (.A_N(_10451_),
    .B(_10452_),
    .C(_10454_),
    .Y(_10455_));
 sky130_fd_sc_hd__nand2_1 _32802_ (.A(_10151_),
    .B(_10152_),
    .Y(_10456_));
 sky130_fd_sc_hd__a21oi_2 _32803_ (.A1(_10156_),
    .A2(_10456_),
    .B1(_10153_),
    .Y(_10457_));
 sky130_fd_sc_hd__buf_4 _32804_ (.A(_19861_),
    .X(_10458_));
 sky130_fd_sc_hd__buf_6 _32805_ (.A(_09972_),
    .X(_10459_));
 sky130_fd_sc_hd__a22oi_4 _32806_ (.A1(_05587_),
    .A2(_10458_),
    .B1(_05589_),
    .B2(_10459_),
    .Y(_10460_));
 sky130_vsdinv _32807_ (.A(_10452_),
    .Y(_10461_));
 sky130_fd_sc_hd__o21ai_2 _32808_ (.A1(_10460_),
    .A2(_10451_),
    .B1(_10461_),
    .Y(_10462_));
 sky130_fd_sc_hd__nand3_4 _32809_ (.A(_10455_),
    .B(_10457_),
    .C(_10462_),
    .Y(_10463_));
 sky130_fd_sc_hd__a21o_1 _32810_ (.A1(_10156_),
    .A2(_10456_),
    .B1(_10153_),
    .X(_10464_));
 sky130_fd_sc_hd__o21ai_2 _32811_ (.A1(_10460_),
    .A2(_10451_),
    .B1(_10452_),
    .Y(_10465_));
 sky130_fd_sc_hd__buf_6 _32812_ (.A(_10449_),
    .X(_10466_));
 sky130_fd_sc_hd__o211ai_4 _32813_ (.A1(_10466_),
    .A2(_10450_),
    .B1(_10461_),
    .C1(_10454_),
    .Y(_10467_));
 sky130_fd_sc_hd__nand3_4 _32814_ (.A(_10464_),
    .B(_10465_),
    .C(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__o21a_1 _32815_ (.A1(_09974_),
    .A2(_09971_),
    .B1(_09977_),
    .X(_10469_));
 sky130_fd_sc_hd__a21o_2 _32816_ (.A1(_10463_),
    .A2(_10468_),
    .B1(_10469_),
    .X(_10470_));
 sky130_fd_sc_hd__nand3_4 _32817_ (.A(_10463_),
    .B(_10468_),
    .C(_10469_),
    .Y(_10471_));
 sky130_fd_sc_hd__nand2_1 _32818_ (.A(_10158_),
    .B(_10147_),
    .Y(_10472_));
 sky130_fd_sc_hd__nand2_4 _32819_ (.A(_10472_),
    .B(_10145_),
    .Y(_10473_));
 sky130_fd_sc_hd__a21oi_4 _32820_ (.A1(_10470_),
    .A2(_10471_),
    .B1(_10473_),
    .Y(_10474_));
 sky130_vsdinv _32821_ (.A(_10468_),
    .Y(_10475_));
 sky130_fd_sc_hd__nand2_1 _32822_ (.A(_10463_),
    .B(_10469_),
    .Y(_10476_));
 sky130_fd_sc_hd__o211a_1 _32823_ (.A1(_10475_),
    .A2(_10476_),
    .B1(_10470_),
    .C1(_10473_),
    .X(_10477_));
 sky130_fd_sc_hd__o22ai_4 _32824_ (.A1(_10447_),
    .A2(_10448_),
    .B1(_10474_),
    .B2(_10477_),
    .Y(_10478_));
 sky130_fd_sc_hd__and2_1 _32825_ (.A(_09991_),
    .B(_09983_),
    .X(_10479_));
 sky130_fd_sc_hd__a21o_1 _32826_ (.A1(_10470_),
    .A2(_10471_),
    .B1(_10473_),
    .X(_10480_));
 sky130_fd_sc_hd__nand3_4 _32827_ (.A(_10473_),
    .B(_10470_),
    .C(_10471_),
    .Y(_10481_));
 sky130_fd_sc_hd__nand3b_4 _32828_ (.A_N(_10479_),
    .B(_10480_),
    .C(_10481_),
    .Y(_10482_));
 sky130_fd_sc_hd__a22oi_4 _32829_ (.A1(_09996_),
    .A2(_10446_),
    .B1(_10478_),
    .B2(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__nor2_1 _32830_ (.A(_10445_),
    .B(_09989_),
    .Y(_10484_));
 sky130_fd_sc_hd__o211a_4 _32831_ (.A1(_09992_),
    .A2(_10484_),
    .B1(_10482_),
    .C1(_10478_),
    .X(_10485_));
 sky130_fd_sc_hd__a21bo_1 _32832_ (.A1(_09956_),
    .A2(_09941_),
    .B1_N(_09945_),
    .X(_10486_));
 sky130_fd_sc_hd__buf_4 _32833_ (.A(\pcpi_mul.rs1[29] ),
    .X(_10487_));
 sky130_fd_sc_hd__buf_4 _32834_ (.A(\pcpi_mul.rs1[28] ),
    .X(_10488_));
 sky130_fd_sc_hd__nand2_1 _32835_ (.A(_05233_),
    .B(_10488_),
    .Y(_10489_));
 sky130_fd_sc_hd__a21o_1 _32836_ (.A1(_19683_),
    .A2(_10487_),
    .B1(_10489_),
    .X(_10490_));
 sky130_fd_sc_hd__nand2_1 _32837_ (.A(_05163_),
    .B(_19834_),
    .Y(_10491_));
 sky130_fd_sc_hd__a21o_1 _32838_ (.A1(_06281_),
    .A2(_19839_),
    .B1(_10491_),
    .X(_10492_));
 sky130_fd_sc_hd__buf_4 _32839_ (.A(_09817_),
    .X(_10493_));
 sky130_fd_sc_hd__nand2_1 _32840_ (.A(_05807_),
    .B(_10493_),
    .Y(_10494_));
 sky130_fd_sc_hd__a21oi_4 _32841_ (.A1(_10490_),
    .A2(_10492_),
    .B1(_10494_),
    .Y(_10495_));
 sky130_vsdinv _32842_ (.A(_09947_),
    .Y(_10496_));
 sky130_fd_sc_hd__clkbuf_8 _32843_ (.A(_10496_),
    .X(_10497_));
 sky130_fd_sc_hd__o211a_2 _32844_ (.A1(_05491_),
    .A2(_10497_),
    .B1(_10490_),
    .C1(_10492_),
    .X(_10498_));
 sky130_fd_sc_hd__nor2_8 _32845_ (.A(_10495_),
    .B(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__nand2_2 _32846_ (.A(_05197_),
    .B(_08787_),
    .Y(_10500_));
 sky130_fd_sc_hd__nand2_2 _32847_ (.A(_05562_),
    .B(_09358_),
    .Y(_10501_));
 sky130_fd_sc_hd__nor2_4 _32848_ (.A(_10500_),
    .B(_10501_),
    .Y(_10502_));
 sky130_fd_sc_hd__and2_1 _32849_ (.A(_10500_),
    .B(_10501_),
    .X(_10503_));
 sky130_fd_sc_hd__buf_6 _32850_ (.A(\pcpi_mul.rs1[30] ),
    .X(_10504_));
 sky130_fd_sc_hd__nand2_2 _32851_ (.A(net476),
    .B(_10504_),
    .Y(_10505_));
 sky130_vsdinv _32852_ (.A(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__o21ai_2 _32853_ (.A1(_10502_),
    .A2(_10503_),
    .B1(_10506_),
    .Y(_10507_));
 sky130_fd_sc_hd__or2_2 _32854_ (.A(_10500_),
    .B(_10501_),
    .X(_10508_));
 sky130_fd_sc_hd__nand2_2 _32855_ (.A(_10500_),
    .B(_10501_),
    .Y(_10509_));
 sky130_fd_sc_hd__nand3_2 _32856_ (.A(_10508_),
    .B(_10505_),
    .C(_10509_),
    .Y(_10510_));
 sky130_fd_sc_hd__a21oi_2 _32857_ (.A1(_09939_),
    .A2(_09935_),
    .B1(_09937_),
    .Y(_10511_));
 sky130_fd_sc_hd__nand3_4 _32858_ (.A(_10507_),
    .B(_10510_),
    .C(_10511_),
    .Y(_10512_));
 sky130_fd_sc_hd__o21ai_2 _32859_ (.A1(_10502_),
    .A2(_10503_),
    .B1(_10505_),
    .Y(_10513_));
 sky130_fd_sc_hd__nand3_2 _32860_ (.A(_10508_),
    .B(_10506_),
    .C(_10509_),
    .Y(_10514_));
 sky130_fd_sc_hd__a21o_1 _32861_ (.A1(_09939_),
    .A2(_09935_),
    .B1(_09937_),
    .X(_10515_));
 sky130_fd_sc_hd__nand3_4 _32862_ (.A(_10513_),
    .B(_10514_),
    .C(_10515_),
    .Y(_10516_));
 sky130_fd_sc_hd__nand3_4 _32863_ (.A(_10499_),
    .B(_10512_),
    .C(_10516_),
    .Y(_10517_));
 sky130_fd_sc_hd__a21o_2 _32864_ (.A1(_10516_),
    .A2(_10512_),
    .B1(_10499_),
    .X(_10518_));
 sky130_fd_sc_hd__nand3_4 _32865_ (.A(_10486_),
    .B(_10517_),
    .C(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__nand2_2 _32866_ (.A(_10518_),
    .B(_10517_),
    .Y(_10520_));
 sky130_fd_sc_hd__a21boi_4 _32867_ (.A1(_09956_),
    .A2(_09941_),
    .B1_N(_09945_),
    .Y(_10521_));
 sky130_fd_sc_hd__o21bai_4 _32868_ (.A1(_09948_),
    .A2(_09951_),
    .B1_N(_09954_),
    .Y(_10522_));
 sky130_fd_sc_hd__a21boi_4 _32869_ (.A1(_10520_),
    .A2(_10521_),
    .B1_N(_10522_),
    .Y(_10523_));
 sky130_fd_sc_hd__nand2_1 _32870_ (.A(_10520_),
    .B(_10521_),
    .Y(_10524_));
 sky130_fd_sc_hd__a21oi_2 _32871_ (.A1(_10524_),
    .A2(_10519_),
    .B1(_10522_),
    .Y(_10525_));
 sky130_fd_sc_hd__a21oi_2 _32872_ (.A1(_10519_),
    .A2(_10523_),
    .B1(_10525_),
    .Y(_10526_));
 sky130_fd_sc_hd__o21ai_2 _32873_ (.A1(_10483_),
    .A2(_10485_),
    .B1(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__a21oi_2 _32874_ (.A1(_10172_),
    .A2(_10179_),
    .B1(_10184_),
    .Y(_10528_));
 sky130_fd_sc_hd__o21ai_2 _32875_ (.A1(_10445_),
    .A2(_09989_),
    .B1(_09997_),
    .Y(_10529_));
 sky130_fd_sc_hd__a21o_1 _32876_ (.A1(_10478_),
    .A2(_10482_),
    .B1(_10529_),
    .X(_10530_));
 sky130_fd_sc_hd__a21o_1 _32877_ (.A1(_10524_),
    .A2(_10519_),
    .B1(_10522_),
    .X(_10531_));
 sky130_fd_sc_hd__nand2_1 _32878_ (.A(_10523_),
    .B(_10519_),
    .Y(_10532_));
 sky130_fd_sc_hd__nand2_4 _32879_ (.A(_10531_),
    .B(_10532_),
    .Y(_10533_));
 sky130_fd_sc_hd__nand3_4 _32880_ (.A(_10478_),
    .B(_10482_),
    .C(_10529_),
    .Y(_10534_));
 sky130_fd_sc_hd__nand3_2 _32881_ (.A(_10530_),
    .B(_10533_),
    .C(_10534_),
    .Y(_10535_));
 sky130_fd_sc_hd__nand3_4 _32882_ (.A(_10527_),
    .B(_10528_),
    .C(_10535_),
    .Y(_10536_));
 sky130_fd_sc_hd__and3_1 _32883_ (.A(_10524_),
    .B(_10519_),
    .C(_10522_),
    .X(_10537_));
 sky130_fd_sc_hd__o22ai_2 _32884_ (.A1(_10537_),
    .A2(_10525_),
    .B1(_10483_),
    .B2(_10485_),
    .Y(_10538_));
 sky130_fd_sc_hd__nand2_1 _32885_ (.A(_10185_),
    .B(_10178_),
    .Y(_10539_));
 sky130_fd_sc_hd__nand3_2 _32886_ (.A(_10530_),
    .B(_10526_),
    .C(_10534_),
    .Y(_10540_));
 sky130_fd_sc_hd__nand3_2 _32887_ (.A(_10538_),
    .B(_10539_),
    .C(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__nand2_1 _32888_ (.A(_10536_),
    .B(_10541_),
    .Y(_10542_));
 sky130_fd_sc_hd__nand2_4 _32889_ (.A(_10011_),
    .B(_10010_),
    .Y(_10543_));
 sky130_vsdinv _32890_ (.A(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__nand2_4 _32891_ (.A(_10542_),
    .B(_10544_),
    .Y(_10545_));
 sky130_fd_sc_hd__buf_2 _32892_ (.A(_10541_),
    .X(_10546_));
 sky130_fd_sc_hd__nand3_4 _32893_ (.A(_10536_),
    .B(_10546_),
    .C(_10543_),
    .Y(_10547_));
 sky130_fd_sc_hd__nand2_1 _32894_ (.A(_10545_),
    .B(_10547_),
    .Y(_10548_));
 sky130_fd_sc_hd__nand2_2 _32895_ (.A(_10444_),
    .B(_10548_),
    .Y(_10549_));
 sky130_vsdinv _32896_ (.A(_10546_),
    .Y(_10550_));
 sky130_fd_sc_hd__nand2_2 _32897_ (.A(_10536_),
    .B(_10543_),
    .Y(_10551_));
 sky130_fd_sc_hd__o2111ai_4 _32898_ (.A1(_10550_),
    .A2(_10551_),
    .B1(_10443_),
    .C1(_10432_),
    .D1(_10545_),
    .Y(_10552_));
 sky130_fd_sc_hd__nand3_4 _32899_ (.A(_10247_),
    .B(_10549_),
    .C(_10552_),
    .Y(_10553_));
 sky130_fd_sc_hd__nand3_2 _32900_ (.A(_10444_),
    .B(_10545_),
    .C(_10547_),
    .Y(_10554_));
 sky130_fd_sc_hd__a21oi_2 _32901_ (.A1(_10192_),
    .A2(_10195_),
    .B1(_10197_),
    .Y(_10555_));
 sky130_fd_sc_hd__a31oi_4 _32902_ (.A1(_10018_),
    .A2(_10198_),
    .A3(_10022_),
    .B1(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__a21oi_2 _32903_ (.A1(_10536_),
    .A2(_10546_),
    .B1(_10543_),
    .Y(_10557_));
 sky130_fd_sc_hd__and3_1 _32904_ (.A(_10005_),
    .B(_10009_),
    .C(_10010_),
    .X(_10558_));
 sky130_fd_sc_hd__o211a_1 _32905_ (.A1(_10003_),
    .A2(_10558_),
    .B1(_10546_),
    .C1(_10536_),
    .X(_10559_));
 sky130_fd_sc_hd__o211ai_4 _32906_ (.A1(_10557_),
    .A2(_10559_),
    .B1(_10432_),
    .C1(_10443_),
    .Y(_10560_));
 sky130_fd_sc_hd__nand3_4 _32907_ (.A(_10554_),
    .B(_10556_),
    .C(_10560_),
    .Y(_10561_));
 sky130_fd_sc_hd__nand2_4 _32908_ (.A(_09965_),
    .B(_09961_),
    .Y(_10562_));
 sky130_fd_sc_hd__nand2_4 _32909_ (.A(_10209_),
    .B(_10021_),
    .Y(_10563_));
 sky130_fd_sc_hd__xor2_4 _32910_ (.A(_10562_),
    .B(_10563_),
    .X(_10564_));
 sky130_fd_sc_hd__nand3_2 _32911_ (.A(_10553_),
    .B(_10561_),
    .C(_10564_),
    .Y(_10565_));
 sky130_vsdinv _32912_ (.A(_10562_),
    .Y(_10566_));
 sky130_vsdinv _32913_ (.A(_10563_),
    .Y(_10567_));
 sky130_fd_sc_hd__nor2_4 _32914_ (.A(_10566_),
    .B(_10567_),
    .Y(_10568_));
 sky130_fd_sc_hd__nor2_1 _32915_ (.A(_10562_),
    .B(_10563_),
    .Y(_10569_));
 sky130_fd_sc_hd__o2bb2ai_2 _32916_ (.A1_N(_10553_),
    .A2_N(_10561_),
    .B1(_10568_),
    .B2(_10569_),
    .Y(_10570_));
 sky130_fd_sc_hd__o211ai_4 _32917_ (.A1(_10244_),
    .A2(_10245_),
    .B1(_10565_),
    .C1(_10570_),
    .Y(_10571_));
 sky130_fd_sc_hd__a21oi_2 _32918_ (.A1(_10219_),
    .A2(_10203_),
    .B1(_10244_),
    .Y(_10572_));
 sky130_fd_sc_hd__nor2_1 _32919_ (.A(_10562_),
    .B(_10567_),
    .Y(_10573_));
 sky130_fd_sc_hd__nor2_1 _32920_ (.A(_10566_),
    .B(_10563_),
    .Y(_10574_));
 sky130_fd_sc_hd__o2bb2ai_2 _32921_ (.A1_N(_10553_),
    .A2_N(_10561_),
    .B1(_10573_),
    .B2(_10574_),
    .Y(_10575_));
 sky130_fd_sc_hd__nand3b_2 _32922_ (.A_N(_10564_),
    .B(_10553_),
    .C(_10561_),
    .Y(_10576_));
 sky130_fd_sc_hd__nand3_4 _32923_ (.A(_10572_),
    .B(_10575_),
    .C(_10576_),
    .Y(_10577_));
 sky130_fd_sc_hd__o2bb2ai_4 _32924_ (.A1_N(_10571_),
    .A2_N(_10577_),
    .B1(_10213_),
    .B2(_10215_),
    .Y(_10578_));
 sky130_fd_sc_hd__nand3_4 _32925_ (.A(_10577_),
    .B(_10571_),
    .C(_10224_),
    .Y(_10579_));
 sky130_fd_sc_hd__nand2_1 _32926_ (.A(_10223_),
    .B(_09896_),
    .Y(_10580_));
 sky130_fd_sc_hd__nand2_2 _32927_ (.A(_10580_),
    .B(_10231_),
    .Y(_10581_));
 sky130_fd_sc_hd__a21oi_2 _32928_ (.A1(_10578_),
    .A2(_10579_),
    .B1(_10581_),
    .Y(_10582_));
 sky130_vsdinv _32929_ (.A(_10231_),
    .Y(_10583_));
 sky130_fd_sc_hd__o211a_1 _32930_ (.A1(_10583_),
    .A2(_10235_),
    .B1(_10579_),
    .C1(_10578_),
    .X(_10584_));
 sky130_fd_sc_hd__nor2_4 _32931_ (.A(_10582_),
    .B(_10584_),
    .Y(_10585_));
 sky130_fd_sc_hd__nor2_2 _32932_ (.A(_09575_),
    .B(_09909_),
    .Y(_10586_));
 sky130_fd_sc_hd__o2bb2ai_2 _32933_ (.A1_N(_09575_),
    .A2_N(_09909_),
    .B1(_09912_),
    .B2(_09914_),
    .Y(_10587_));
 sky130_fd_sc_hd__o2111ai_4 _32934_ (.A1(_10586_),
    .A2(_10587_),
    .B1(_09917_),
    .C1(_10240_),
    .D1(_10237_),
    .Y(_10588_));
 sky130_fd_sc_hd__a21bo_1 _32935_ (.A1(_09915_),
    .A2(_10237_),
    .B1_N(_10240_),
    .X(_10589_));
 sky130_fd_sc_hd__o21ai_1 _32936_ (.A1(_10588_),
    .A2(_09925_),
    .B1(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__nor2_1 _32937_ (.A(_10585_),
    .B(_10590_),
    .Y(_10591_));
 sky130_fd_sc_hd__and2_1 _32938_ (.A(_10590_),
    .B(_10585_),
    .X(_10592_));
 sky130_fd_sc_hd__nor2_2 _32939_ (.A(_10591_),
    .B(_10592_),
    .Y(_02649_));
 sky130_vsdinv _32940_ (.A(_10424_),
    .Y(_10593_));
 sky130_fd_sc_hd__a21bo_1 _32941_ (.A1(_10512_),
    .A2(_10499_),
    .B1_N(_10516_),
    .X(_10594_));
 sky130_fd_sc_hd__and4_1 _32942_ (.A(_05117_),
    .B(_05119_),
    .C(_10504_),
    .D(_19834_),
    .X(_10595_));
 sky130_vsdinv _32943_ (.A(\pcpi_mul.rs1[30] ),
    .Y(_10596_));
 sky130_fd_sc_hd__buf_6 _32944_ (.A(_10596_),
    .X(_10597_));
 sky130_fd_sc_hd__clkbuf_4 _32945_ (.A(\pcpi_mul.rs1[29] ),
    .X(_10598_));
 sky130_fd_sc_hd__nand2_1 _32946_ (.A(_06281_),
    .B(_10598_),
    .Y(_10599_));
 sky130_fd_sc_hd__o21a_1 _32947_ (.A1(_05153_),
    .A2(_10597_),
    .B1(_10599_),
    .X(_10600_));
 sky130_fd_sc_hd__buf_4 _32948_ (.A(_19838_),
    .X(_10601_));
 sky130_fd_sc_hd__nand2_1 _32949_ (.A(_05807_),
    .B(_10601_),
    .Y(_10602_));
 sky130_vsdinv _32950_ (.A(_10602_),
    .Y(_10603_));
 sky130_fd_sc_hd__o21ai_1 _32951_ (.A1(_10595_),
    .A2(_10600_),
    .B1(_10603_),
    .Y(_10604_));
 sky130_fd_sc_hd__o21ai_1 _32952_ (.A1(_05153_),
    .A2(_10597_),
    .B1(_10599_),
    .Y(_10605_));
 sky130_fd_sc_hd__nand3b_2 _32953_ (.A_N(_10595_),
    .B(_10602_),
    .C(_10605_),
    .Y(_10606_));
 sky130_fd_sc_hd__nand2_2 _32954_ (.A(_10604_),
    .B(_10606_),
    .Y(_10607_));
 sky130_fd_sc_hd__a21oi_4 _32955_ (.A1(_10506_),
    .A2(_10509_),
    .B1(_10502_),
    .Y(_10608_));
 sky130_fd_sc_hd__nand2_2 _32956_ (.A(_19670_),
    .B(_09358_),
    .Y(_10609_));
 sky130_fd_sc_hd__nand2_2 _32957_ (.A(_05358_),
    .B(_09947_),
    .Y(_10610_));
 sky130_fd_sc_hd__or2_2 _32958_ (.A(_10609_),
    .B(_10610_),
    .X(_10611_));
 sky130_fd_sc_hd__nand2_4 _32959_ (.A(_10609_),
    .B(_10610_),
    .Y(_10612_));
 sky130_fd_sc_hd__buf_4 _32960_ (.A(\pcpi_mul.rs1[31] ),
    .X(_10613_));
 sky130_fd_sc_hd__nand2_1 _32961_ (.A(net476),
    .B(_10613_),
    .Y(_10614_));
 sky130_vsdinv _32962_ (.A(_10614_),
    .Y(_10615_));
 sky130_fd_sc_hd__nand3_2 _32963_ (.A(_10611_),
    .B(_10612_),
    .C(_10615_),
    .Y(_10616_));
 sky130_vsdinv _32964_ (.A(_19847_),
    .Y(_10617_));
 sky130_fd_sc_hd__nand3_4 _32965_ (.A(_05791_),
    .B(_05792_),
    .C(_09817_),
    .Y(_10618_));
 sky130_fd_sc_hd__o21ai_1 _32966_ (.A1(_10617_),
    .A2(_10618_),
    .B1(_10612_),
    .Y(_10619_));
 sky130_fd_sc_hd__nand2_1 _32967_ (.A(_10619_),
    .B(_10614_),
    .Y(_10620_));
 sky130_fd_sc_hd__nand3b_4 _32968_ (.A_N(_10608_),
    .B(_10616_),
    .C(_10620_),
    .Y(_10621_));
 sky130_fd_sc_hd__nand3_2 _32969_ (.A(_10611_),
    .B(_10612_),
    .C(_10614_),
    .Y(_10622_));
 sky130_fd_sc_hd__nand2_1 _32970_ (.A(_10619_),
    .B(_10615_),
    .Y(_10623_));
 sky130_fd_sc_hd__nand3_4 _32971_ (.A(_10622_),
    .B(_10623_),
    .C(_10608_),
    .Y(_10624_));
 sky130_fd_sc_hd__nand3_2 _32972_ (.A(_10607_),
    .B(_10621_),
    .C(_10624_),
    .Y(_10625_));
 sky130_fd_sc_hd__nand2_1 _32973_ (.A(_10621_),
    .B(_10624_),
    .Y(_10626_));
 sky130_fd_sc_hd__and2_1 _32974_ (.A(_10604_),
    .B(_10606_),
    .X(_10627_));
 sky130_fd_sc_hd__nand2_1 _32975_ (.A(_10626_),
    .B(_10627_),
    .Y(_10628_));
 sky130_fd_sc_hd__nand3_4 _32976_ (.A(_10594_),
    .B(_10625_),
    .C(_10628_),
    .Y(_10629_));
 sky130_fd_sc_hd__nand2_1 _32977_ (.A(_10626_),
    .B(_10607_),
    .Y(_10630_));
 sky130_fd_sc_hd__a21boi_4 _32978_ (.A1(_10499_),
    .A2(_10512_),
    .B1_N(_10516_),
    .Y(_10631_));
 sky130_fd_sc_hd__nand3_2 _32979_ (.A(_10627_),
    .B(_10621_),
    .C(_10624_),
    .Y(_10632_));
 sky130_fd_sc_hd__nand3_4 _32980_ (.A(_10630_),
    .B(_10631_),
    .C(_10632_),
    .Y(_10633_));
 sky130_fd_sc_hd__nor2_1 _32981_ (.A(_10489_),
    .B(_10491_),
    .Y(_10634_));
 sky130_fd_sc_hd__nor2_1 _32982_ (.A(_10634_),
    .B(_10495_),
    .Y(_10635_));
 sky130_fd_sc_hd__a21boi_4 _32983_ (.A1(_10629_),
    .A2(_10633_),
    .B1_N(_10635_),
    .Y(_10636_));
 sky130_vsdinv _32984_ (.A(_10636_),
    .Y(_10637_));
 sky130_fd_sc_hd__o21a_1 _32985_ (.A1(_10634_),
    .A2(_10495_),
    .B1(_10633_),
    .X(_10638_));
 sky130_fd_sc_hd__nand2_2 _32986_ (.A(_10638_),
    .B(_10629_),
    .Y(_10639_));
 sky130_fd_sc_hd__nand3_4 _32987_ (.A(_05440_),
    .B(_19664_),
    .C(_09972_),
    .Y(_10640_));
 sky130_fd_sc_hd__nor2_8 _32988_ (.A(_09806_),
    .B(_10640_),
    .Y(_10641_));
 sky130_fd_sc_hd__nand2_2 _32989_ (.A(_19667_),
    .B(_09079_),
    .Y(_10642_));
 sky130_fd_sc_hd__buf_4 _32990_ (.A(_09076_),
    .X(_10643_));
 sky130_fd_sc_hd__a22o_1 _32991_ (.A1(_05837_),
    .A2(_10453_),
    .B1(_19665_),
    .B2(_10643_),
    .X(_10644_));
 sky130_fd_sc_hd__nand3b_2 _32992_ (.A_N(_10641_),
    .B(_10642_),
    .C(_10644_),
    .Y(_10645_));
 sky130_fd_sc_hd__o22a_1 _32993_ (.A1(_08079_),
    .A2(_10397_),
    .B1(_10399_),
    .B2(_10396_),
    .X(_10646_));
 sky130_fd_sc_hd__a22oi_4 _32994_ (.A1(_06076_),
    .A2(_19858_),
    .B1(_06077_),
    .B2(_19854_),
    .Y(_10647_));
 sky130_vsdinv _32995_ (.A(_10642_),
    .Y(_10648_));
 sky130_fd_sc_hd__o21ai_2 _32996_ (.A1(_10647_),
    .A2(_10641_),
    .B1(_10648_),
    .Y(_10649_));
 sky130_fd_sc_hd__nand3_4 _32997_ (.A(_10645_),
    .B(_10646_),
    .C(_10649_),
    .Y(_10650_));
 sky130_fd_sc_hd__o21ai_2 _32998_ (.A1(_10647_),
    .A2(_10641_),
    .B1(_10642_),
    .Y(_10651_));
 sky130_fd_sc_hd__buf_6 _32999_ (.A(_09806_),
    .X(_10652_));
 sky130_fd_sc_hd__o211ai_4 _33000_ (.A1(_10652_),
    .A2(_10640_),
    .B1(_10648_),
    .C1(_10644_),
    .Y(_10653_));
 sky130_fd_sc_hd__buf_4 _33001_ (.A(_08079_),
    .X(_10654_));
 sky130_fd_sc_hd__o22ai_4 _33002_ (.A1(_10654_),
    .A2(_10397_),
    .B1(_10399_),
    .B2(_10396_),
    .Y(_10655_));
 sky130_fd_sc_hd__nand3_4 _33003_ (.A(_10651_),
    .B(_10653_),
    .C(_10655_),
    .Y(_10656_));
 sky130_fd_sc_hd__nand2_1 _33004_ (.A(_10650_),
    .B(_10656_),
    .Y(_10657_));
 sky130_fd_sc_hd__a21oi_4 _33005_ (.A1(_10454_),
    .A2(_10461_),
    .B1(_10451_),
    .Y(_10658_));
 sky130_fd_sc_hd__nand2_4 _33006_ (.A(_10657_),
    .B(_10658_),
    .Y(_10659_));
 sky130_vsdinv _33007_ (.A(_10658_),
    .Y(_10660_));
 sky130_fd_sc_hd__nand3_4 _33008_ (.A(_10650_),
    .B(_10656_),
    .C(_10660_),
    .Y(_10661_));
 sky130_fd_sc_hd__nand2_4 _33009_ (.A(_10659_),
    .B(_10661_),
    .Y(_10662_));
 sky130_fd_sc_hd__a21o_1 _33010_ (.A1(_10139_),
    .A2(_10142_),
    .B1(_10137_),
    .X(_10663_));
 sky130_fd_sc_hd__o31a_1 _33011_ (.A1(_10387_),
    .A2(_10385_),
    .A3(_10386_),
    .B1(_10663_),
    .X(_10664_));
 sky130_fd_sc_hd__o21ai_2 _33012_ (.A1(_10385_),
    .A2(_10386_),
    .B1(_10387_),
    .Y(_10665_));
 sky130_fd_sc_hd__a22oi_4 _33013_ (.A1(_10664_),
    .A2(_10665_),
    .B1(_10392_),
    .B2(_10406_),
    .Y(_10666_));
 sky130_fd_sc_hd__nand2_1 _33014_ (.A(_10662_),
    .B(_10666_),
    .Y(_10667_));
 sky130_fd_sc_hd__nand2_1 _33015_ (.A(_10406_),
    .B(_10392_),
    .Y(_10668_));
 sky130_fd_sc_hd__nand2_2 _33016_ (.A(_10668_),
    .B(_10393_),
    .Y(_10669_));
 sky130_fd_sc_hd__nand3_4 _33017_ (.A(_10669_),
    .B(_10661_),
    .C(_10659_),
    .Y(_10670_));
 sky130_fd_sc_hd__nand2_1 _33018_ (.A(_10476_),
    .B(_10468_),
    .Y(_10671_));
 sky130_fd_sc_hd__a21oi_2 _33019_ (.A1(_10667_),
    .A2(_10670_),
    .B1(_10671_),
    .Y(_10672_));
 sky130_vsdinv _33020_ (.A(_10671_),
    .Y(_10673_));
 sky130_fd_sc_hd__a21oi_4 _33021_ (.A1(_10659_),
    .A2(_10661_),
    .B1(_10669_),
    .Y(_10674_));
 sky130_fd_sc_hd__nor2_8 _33022_ (.A(_10666_),
    .B(_10662_),
    .Y(_10675_));
 sky130_fd_sc_hd__nor3_4 _33023_ (.A(_10673_),
    .B(_10674_),
    .C(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__o21ai_4 _33024_ (.A1(_10479_),
    .A2(_10474_),
    .B1(_10481_),
    .Y(_10677_));
 sky130_fd_sc_hd__o21bai_4 _33025_ (.A1(_10672_),
    .A2(_10676_),
    .B1_N(_10677_),
    .Y(_10678_));
 sky130_fd_sc_hd__o21ai_2 _33026_ (.A1(_10674_),
    .A2(_10675_),
    .B1(_10673_),
    .Y(_10679_));
 sky130_fd_sc_hd__a21oi_4 _33027_ (.A1(_10662_),
    .A2(_10666_),
    .B1(_10673_),
    .Y(_10680_));
 sky130_fd_sc_hd__nand2_2 _33028_ (.A(_10680_),
    .B(_10670_),
    .Y(_10681_));
 sky130_fd_sc_hd__nand3_4 _33029_ (.A(_10679_),
    .B(_10681_),
    .C(_10677_),
    .Y(_10682_));
 sky130_fd_sc_hd__a22oi_4 _33030_ (.A1(_10637_),
    .A2(_10639_),
    .B1(_10678_),
    .B2(_10682_),
    .Y(_10683_));
 sky130_fd_sc_hd__a21oi_2 _33031_ (.A1(_10679_),
    .A2(_10681_),
    .B1(_10677_),
    .Y(_10684_));
 sky130_fd_sc_hd__a21oi_4 _33032_ (.A1(_10629_),
    .A2(_10638_),
    .B1(_10636_),
    .Y(_10685_));
 sky130_fd_sc_hd__nand2_1 _33033_ (.A(_10685_),
    .B(_10682_),
    .Y(_10686_));
 sky130_fd_sc_hd__nor2_2 _33034_ (.A(_10684_),
    .B(_10686_),
    .Y(_10687_));
 sky130_fd_sc_hd__o22ai_4 _33035_ (.A1(_10423_),
    .A2(_10593_),
    .B1(_10683_),
    .B2(_10687_),
    .Y(_10688_));
 sky130_vsdinv _33036_ (.A(_10639_),
    .Y(_10689_));
 sky130_fd_sc_hd__o2bb2ai_4 _33037_ (.A1_N(_10682_),
    .A2_N(_10678_),
    .B1(_10636_),
    .B2(_10689_),
    .Y(_10690_));
 sky130_fd_sc_hd__o21ai_4 _33038_ (.A1(_10421_),
    .A2(_10423_),
    .B1(_10419_),
    .Y(_10691_));
 sky130_fd_sc_hd__nand3_4 _33039_ (.A(_10678_),
    .B(_10685_),
    .C(_10682_),
    .Y(_10692_));
 sky130_fd_sc_hd__nand3_4 _33040_ (.A(_10690_),
    .B(_10691_),
    .C(_10692_),
    .Y(_10693_));
 sky130_fd_sc_hd__nor2_8 _33041_ (.A(_10483_),
    .B(_10533_),
    .Y(_10694_));
 sky130_fd_sc_hd__nor2_8 _33042_ (.A(_10485_),
    .B(_10694_),
    .Y(_10695_));
 sky130_fd_sc_hd__a21oi_2 _33043_ (.A1(_10688_),
    .A2(_10693_),
    .B1(_10695_),
    .Y(_10696_));
 sky130_fd_sc_hd__a21oi_4 _33044_ (.A1(_10690_),
    .A2(_10692_),
    .B1(_10691_),
    .Y(_10697_));
 sky130_fd_sc_hd__nand2_4 _33045_ (.A(_10693_),
    .B(_10695_),
    .Y(_10698_));
 sky130_fd_sc_hd__nor2_2 _33046_ (.A(_10697_),
    .B(_10698_),
    .Y(_10699_));
 sky130_fd_sc_hd__nand3_4 _33047_ (.A(_19631_),
    .B(_07428_),
    .C(_07322_),
    .Y(_10700_));
 sky130_fd_sc_hd__a22o_2 _33048_ (.A1(_07744_),
    .A2(_07330_),
    .B1(_06921_),
    .B2(_07059_),
    .X(_10701_));
 sky130_fd_sc_hd__o21ai_2 _33049_ (.A1(_06810_),
    .A2(_10700_),
    .B1(_10701_),
    .Y(_10702_));
 sky130_fd_sc_hd__nand2_2 _33050_ (.A(_19641_),
    .B(_07052_),
    .Y(_10703_));
 sky130_vsdinv _33051_ (.A(_10703_),
    .Y(_10704_));
 sky130_fd_sc_hd__nand2_4 _33052_ (.A(_10702_),
    .B(_10704_),
    .Y(_10705_));
 sky130_fd_sc_hd__nor2_8 _33053_ (.A(_06809_),
    .B(_10700_),
    .Y(_10706_));
 sky130_fd_sc_hd__nand3b_4 _33054_ (.A_N(_10706_),
    .B(_10703_),
    .C(_10701_),
    .Y(_10707_));
 sky130_fd_sc_hd__a21oi_4 _33055_ (.A1(_10321_),
    .A2(_10323_),
    .B1(_10318_),
    .Y(_10708_));
 sky130_fd_sc_hd__nand3_4 _33056_ (.A(_10705_),
    .B(_10707_),
    .C(_10708_),
    .Y(_10709_));
 sky130_fd_sc_hd__nand2_1 _33057_ (.A(_10702_),
    .B(_10703_),
    .Y(_10710_));
 sky130_fd_sc_hd__nand3b_4 _33058_ (.A_N(_10706_),
    .B(_10704_),
    .C(_10701_),
    .Y(_10711_));
 sky130_fd_sc_hd__nand3b_4 _33059_ (.A_N(_10708_),
    .B(_10710_),
    .C(_10711_),
    .Y(_10712_));
 sky130_fd_sc_hd__nor2_2 _33060_ (.A(_10367_),
    .B(_10359_),
    .Y(_10713_));
 sky130_fd_sc_hd__o2bb2ai_4 _33061_ (.A1_N(_10709_),
    .A2_N(_10712_),
    .B1(_10360_),
    .B2(_10713_),
    .Y(_10714_));
 sky130_fd_sc_hd__a21oi_4 _33062_ (.A1(_10367_),
    .A2(_10368_),
    .B1(_10359_),
    .Y(_10715_));
 sky130_vsdinv _33063_ (.A(_10715_),
    .Y(_10716_));
 sky130_fd_sc_hd__nand3_4 _33064_ (.A(_10712_),
    .B(_10709_),
    .C(_10716_),
    .Y(_10717_));
 sky130_fd_sc_hd__nand2_2 _33065_ (.A(_10381_),
    .B(_10370_),
    .Y(_10718_));
 sky130_fd_sc_hd__a21oi_4 _33066_ (.A1(_10714_),
    .A2(_10717_),
    .B1(_10718_),
    .Y(_10719_));
 sky130_fd_sc_hd__a31oi_4 _33067_ (.A1(_10705_),
    .A2(_10707_),
    .A3(_10708_),
    .B1(_10715_),
    .Y(_10720_));
 sky130_fd_sc_hd__a21oi_1 _33068_ (.A1(_10712_),
    .A2(_10709_),
    .B1(_10716_),
    .Y(_10721_));
 sky130_fd_sc_hd__a221oi_2 _33069_ (.A1(_10720_),
    .A2(_10712_),
    .B1(_10381_),
    .B2(_10370_),
    .C1(_10721_),
    .Y(_10722_));
 sky130_fd_sc_hd__a22oi_4 _33070_ (.A1(_06342_),
    .A2(_07344_),
    .B1(_06618_),
    .B2(_19874_),
    .Y(_10723_));
 sky130_vsdinv _33071_ (.A(_07554_),
    .Y(_10724_));
 sky130_fd_sc_hd__nand3_4 _33072_ (.A(_06896_),
    .B(_06898_),
    .C(_08734_),
    .Y(_10725_));
 sky130_fd_sc_hd__nor2_8 _33073_ (.A(_10724_),
    .B(_10725_),
    .Y(_10726_));
 sky130_fd_sc_hd__nand2_2 _33074_ (.A(_06349_),
    .B(_08062_),
    .Y(_10727_));
 sky130_vsdinv _33075_ (.A(_10727_),
    .Y(_10728_));
 sky130_fd_sc_hd__o21ai_2 _33076_ (.A1(_10723_),
    .A2(_10726_),
    .B1(_10728_),
    .Y(_10729_));
 sky130_vsdinv _33077_ (.A(_10387_),
    .Y(_10730_));
 sky130_fd_sc_hd__a21oi_4 _33078_ (.A1(_10730_),
    .A2(_10389_),
    .B1(_10385_),
    .Y(_10731_));
 sky130_fd_sc_hd__buf_6 _33079_ (.A(_10724_),
    .X(_10732_));
 sky130_fd_sc_hd__buf_4 _33080_ (.A(_07067_),
    .X(_10733_));
 sky130_fd_sc_hd__a22o_2 _33081_ (.A1(_06411_),
    .A2(_07051_),
    .B1(_06169_),
    .B2(_10733_),
    .X(_10734_));
 sky130_fd_sc_hd__o211ai_4 _33082_ (.A1(_10732_),
    .A2(_10725_),
    .B1(_10727_),
    .C1(_10734_),
    .Y(_10735_));
 sky130_fd_sc_hd__nand3_4 _33083_ (.A(_10729_),
    .B(_10731_),
    .C(_10735_),
    .Y(_10736_));
 sky130_fd_sc_hd__buf_4 _33084_ (.A(_07893_),
    .X(_10737_));
 sky130_fd_sc_hd__buf_6 _33085_ (.A(_08056_),
    .X(_10738_));
 sky130_fd_sc_hd__a22oi_4 _33086_ (.A1(_10737_),
    .A2(_19869_),
    .B1(_06336_),
    .B2(_10738_),
    .Y(_10739_));
 sky130_fd_sc_hd__nand2_1 _33087_ (.A(_06883_),
    .B(_10395_),
    .Y(_10740_));
 sky130_fd_sc_hd__nand2_1 _33088_ (.A(_06399_),
    .B(_08336_),
    .Y(_10741_));
 sky130_fd_sc_hd__nor2_2 _33089_ (.A(_10740_),
    .B(_10741_),
    .Y(_10742_));
 sky130_fd_sc_hd__nand2_1 _33090_ (.A(_05732_),
    .B(_19863_),
    .Y(_10743_));
 sky130_fd_sc_hd__o21bai_1 _33091_ (.A1(_10739_),
    .A2(_10742_),
    .B1_N(_10743_),
    .Y(_10744_));
 sky130_fd_sc_hd__buf_4 _33092_ (.A(_08333_),
    .X(_10745_));
 sky130_fd_sc_hd__nand3b_2 _33093_ (.A_N(_10740_),
    .B(_06160_),
    .C(_10745_),
    .Y(_10746_));
 sky130_fd_sc_hd__nand2_2 _33094_ (.A(_10740_),
    .B(_10741_),
    .Y(_10747_));
 sky130_fd_sc_hd__nand3_1 _33095_ (.A(_10746_),
    .B(_10743_),
    .C(_10747_),
    .Y(_10748_));
 sky130_fd_sc_hd__nand2_2 _33096_ (.A(_10744_),
    .B(_10748_),
    .Y(_10749_));
 sky130_fd_sc_hd__nand2_2 _33097_ (.A(_10736_),
    .B(_10749_),
    .Y(_10750_));
 sky130_fd_sc_hd__a21o_1 _33098_ (.A1(_10729_),
    .A2(_10735_),
    .B1(_10731_),
    .X(_10751_));
 sky130_fd_sc_hd__or2b_1 _33099_ (.A(_10750_),
    .B_N(_10751_),
    .X(_10752_));
 sky130_fd_sc_hd__nand2_1 _33100_ (.A(_10751_),
    .B(_10736_),
    .Y(_10753_));
 sky130_vsdinv _33101_ (.A(_10749_),
    .Y(_10754_));
 sky130_fd_sc_hd__nand2_1 _33102_ (.A(_10753_),
    .B(_10754_),
    .Y(_10755_));
 sky130_fd_sc_hd__nand2_2 _33103_ (.A(_10752_),
    .B(_10755_),
    .Y(_10756_));
 sky130_fd_sc_hd__o21ai_2 _33104_ (.A1(_10719_),
    .A2(_10722_),
    .B1(_10756_),
    .Y(_10757_));
 sky130_fd_sc_hd__nand2_4 _33105_ (.A(_10350_),
    .B(_10340_),
    .Y(_10758_));
 sky130_fd_sc_hd__a21o_2 _33106_ (.A1(_10714_),
    .A2(_10717_),
    .B1(_10718_),
    .X(_10759_));
 sky130_fd_sc_hd__nand3_4 _33107_ (.A(_10718_),
    .B(_10714_),
    .C(_10717_),
    .Y(_10760_));
 sky130_fd_sc_hd__nand2_1 _33108_ (.A(_10753_),
    .B(_10749_),
    .Y(_10761_));
 sky130_fd_sc_hd__nand3_2 _33109_ (.A(_10754_),
    .B(_10751_),
    .C(_10736_),
    .Y(_10762_));
 sky130_fd_sc_hd__nand2_2 _33110_ (.A(_10761_),
    .B(_10762_),
    .Y(_10763_));
 sky130_fd_sc_hd__nand3_4 _33111_ (.A(_10759_),
    .B(_10760_),
    .C(_10763_),
    .Y(_10764_));
 sky130_fd_sc_hd__nand3_4 _33112_ (.A(_10757_),
    .B(_10758_),
    .C(_10764_),
    .Y(_10765_));
 sky130_vsdinv _33113_ (.A(_10762_),
    .Y(_10766_));
 sky130_vsdinv _33114_ (.A(_10761_),
    .Y(_10767_));
 sky130_fd_sc_hd__o22ai_4 _33115_ (.A1(_10766_),
    .A2(_10767_),
    .B1(_10719_),
    .B2(_10722_),
    .Y(_10768_));
 sky130_fd_sc_hd__a21oi_4 _33116_ (.A1(_10339_),
    .A2(_10335_),
    .B1(_10334_),
    .Y(_10769_));
 sky130_fd_sc_hd__nand3_2 _33117_ (.A(_10759_),
    .B(_10760_),
    .C(_10756_),
    .Y(_10770_));
 sky130_fd_sc_hd__nand3_4 _33118_ (.A(_10768_),
    .B(_10769_),
    .C(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__nor2_8 _33119_ (.A(_10408_),
    .B(_10413_),
    .Y(_10772_));
 sky130_fd_sc_hd__nor2_8 _33120_ (.A(_10414_),
    .B(_10772_),
    .Y(_10773_));
 sky130_fd_sc_hd__a21oi_2 _33121_ (.A1(_10765_),
    .A2(_10771_),
    .B1(_10773_),
    .Y(_10774_));
 sky130_fd_sc_hd__nand3_4 _33122_ (.A(_10765_),
    .B(_10771_),
    .C(_10773_),
    .Y(_10775_));
 sky130_vsdinv _33123_ (.A(_10775_),
    .Y(_10776_));
 sky130_vsdinv _33124_ (.A(_10314_),
    .Y(_10777_));
 sky130_fd_sc_hd__and3_1 _33125_ (.A(_10310_),
    .B(_10322_),
    .C(_10324_),
    .X(_10778_));
 sky130_fd_sc_hd__nand2_2 _33126_ (.A(_09191_),
    .B(_05660_),
    .Y(_10779_));
 sky130_fd_sc_hd__nand2_2 _33127_ (.A(_09516_),
    .B(_19903_),
    .Y(_10780_));
 sky130_fd_sc_hd__nor2_4 _33128_ (.A(_10779_),
    .B(_10780_),
    .Y(_10781_));
 sky130_fd_sc_hd__nand2_2 _33129_ (.A(_19615_),
    .B(_19900_),
    .Y(_10782_));
 sky130_fd_sc_hd__nand2_4 _33130_ (.A(_10779_),
    .B(_10780_),
    .Y(_10783_));
 sky130_fd_sc_hd__nand3b_2 _33131_ (.A_N(_10781_),
    .B(_10782_),
    .C(_10783_),
    .Y(_10784_));
 sky130_fd_sc_hd__a21oi_2 _33132_ (.A1(_10305_),
    .A2(_10304_),
    .B1(_10302_),
    .Y(_10785_));
 sky130_fd_sc_hd__a22oi_4 _33133_ (.A1(_19607_),
    .A2(_06105_),
    .B1(_07984_),
    .B2(_06264_),
    .Y(_10786_));
 sky130_vsdinv _33134_ (.A(_10782_),
    .Y(_10787_));
 sky130_fd_sc_hd__o21ai_2 _33135_ (.A1(_10786_),
    .A2(_10781_),
    .B1(_10787_),
    .Y(_10788_));
 sky130_fd_sc_hd__nand3_4 _33136_ (.A(_10784_),
    .B(_10785_),
    .C(_10788_),
    .Y(_10789_));
 sky130_fd_sc_hd__nor2_2 _33137_ (.A(_10303_),
    .B(_10308_),
    .Y(_10790_));
 sky130_fd_sc_hd__nand3_4 _33138_ (.A(_09191_),
    .B(_09516_),
    .C(_05801_),
    .Y(_10791_));
 sky130_fd_sc_hd__o211ai_4 _33139_ (.A1(net449),
    .A2(_10791_),
    .B1(_10783_),
    .C1(_10787_),
    .Y(_10792_));
 sky130_fd_sc_hd__o21ai_2 _33140_ (.A1(_10786_),
    .A2(_10781_),
    .B1(_10782_),
    .Y(_10793_));
 sky130_fd_sc_hd__o211ai_4 _33141_ (.A1(_10302_),
    .A2(_10790_),
    .B1(_10792_),
    .C1(_10793_),
    .Y(_10794_));
 sky130_fd_sc_hd__a22oi_4 _33142_ (.A1(_07978_),
    .A2(_19898_),
    .B1(_19625_),
    .B2(_06788_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand2_4 _33143_ (.A(_07822_),
    .B(_06648_),
    .Y(_10796_));
 sky130_fd_sc_hd__nand2_4 _33144_ (.A(_07827_),
    .B(_07502_),
    .Y(_10797_));
 sky130_fd_sc_hd__nor2_8 _33145_ (.A(_10796_),
    .B(_10797_),
    .Y(_10798_));
 sky130_fd_sc_hd__a211o_2 _33146_ (.A1(_19628_),
    .A2(_19892_),
    .B1(_10795_),
    .C1(_10798_),
    .X(_10799_));
 sky130_fd_sc_hd__nor2_8 _33147_ (.A(_07041_),
    .B(net440),
    .Y(_10800_));
 sky130_fd_sc_hd__o21ai_2 _33148_ (.A1(_10795_),
    .A2(_10798_),
    .B1(_10800_),
    .Y(_10801_));
 sky130_fd_sc_hd__nand2_4 _33149_ (.A(_10799_),
    .B(_10801_),
    .Y(_10802_));
 sky130_fd_sc_hd__a21o_2 _33150_ (.A1(_10789_),
    .A2(_10794_),
    .B1(_10802_),
    .X(_10803_));
 sky130_fd_sc_hd__buf_2 _33151_ (.A(_10794_),
    .X(_10804_));
 sky130_fd_sc_hd__nand3_4 _33152_ (.A(_10802_),
    .B(_10789_),
    .C(_10804_),
    .Y(_10805_));
 sky130_fd_sc_hd__nand2_2 _33153_ (.A(_10292_),
    .B(_10264_),
    .Y(_10806_));
 sky130_fd_sc_hd__a21oi_4 _33154_ (.A1(_10803_),
    .A2(_10805_),
    .B1(_10806_),
    .Y(_10807_));
 sky130_fd_sc_hd__o211a_4 _33155_ (.A1(_10293_),
    .A2(_10272_),
    .B1(_10805_),
    .C1(_10803_),
    .X(_10808_));
 sky130_fd_sc_hd__o22ai_4 _33156_ (.A1(_10777_),
    .A2(_10778_),
    .B1(_10807_),
    .B2(_10808_),
    .Y(_10809_));
 sky130_fd_sc_hd__a21oi_2 _33157_ (.A1(_10789_),
    .A2(_10804_),
    .B1(_10802_),
    .Y(_10810_));
 sky130_fd_sc_hd__o21a_1 _33158_ (.A1(_10795_),
    .A2(_10798_),
    .B1(_10800_),
    .X(_10811_));
 sky130_fd_sc_hd__nor3_1 _33159_ (.A(_10795_),
    .B(_10798_),
    .C(_10800_),
    .Y(_10812_));
 sky130_fd_sc_hd__o211a_1 _33160_ (.A1(_10811_),
    .A2(_10812_),
    .B1(_10804_),
    .C1(_10789_),
    .X(_10813_));
 sky130_fd_sc_hd__nor2_2 _33161_ (.A(_10272_),
    .B(_10293_),
    .Y(_10814_));
 sky130_fd_sc_hd__o21ai_4 _33162_ (.A1(_10810_),
    .A2(_10813_),
    .B1(_10814_),
    .Y(_10815_));
 sky130_fd_sc_hd__nand3_4 _33163_ (.A(_10803_),
    .B(_10806_),
    .C(_10805_),
    .Y(_10816_));
 sky130_fd_sc_hd__nand2_1 _33164_ (.A(_10327_),
    .B(_10314_),
    .Y(_10817_));
 sky130_fd_sc_hd__nand2_4 _33165_ (.A(_10817_),
    .B(_10310_),
    .Y(_10818_));
 sky130_fd_sc_hd__nand3_4 _33166_ (.A(_10815_),
    .B(_10816_),
    .C(_10818_),
    .Y(_10819_));
 sky130_fd_sc_hd__nand2_8 _33167_ (.A(_19582_),
    .B(_07828_),
    .Y(_10820_));
 sky130_fd_sc_hd__nand2_8 _33168_ (.A(_19586_),
    .B(_19923_),
    .Y(_10821_));
 sky130_fd_sc_hd__or2_2 _33169_ (.A(_10820_),
    .B(_10821_),
    .X(_10822_));
 sky130_fd_sc_hd__nand2_4 _33170_ (.A(_10820_),
    .B(_10821_),
    .Y(_10823_));
 sky130_fd_sc_hd__nand2_4 _33171_ (.A(_19591_),
    .B(_07008_),
    .Y(_10824_));
 sky130_vsdinv _33172_ (.A(_10824_),
    .Y(_10825_));
 sky130_fd_sc_hd__nand3_2 _33173_ (.A(_10822_),
    .B(_10823_),
    .C(_10825_),
    .Y(_10826_));
 sky130_fd_sc_hd__buf_6 _33174_ (.A(\pcpi_mul.rs2[30] ),
    .X(_10827_));
 sky130_fd_sc_hd__buf_4 _33175_ (.A(_10827_),
    .X(_10828_));
 sky130_fd_sc_hd__a22oi_4 _33176_ (.A1(_19576_),
    .A2(_19933_),
    .B1(_10828_),
    .B2(_07759_),
    .Y(_10829_));
 sky130_fd_sc_hd__clkbuf_4 _33177_ (.A(\pcpi_mul.rs2[31] ),
    .X(_10830_));
 sky130_fd_sc_hd__nand2_2 _33178_ (.A(_10830_),
    .B(_05204_),
    .Y(_10831_));
 sky130_fd_sc_hd__nand2_2 _33179_ (.A(_19579_),
    .B(_05441_),
    .Y(_10832_));
 sky130_fd_sc_hd__nor2_8 _33180_ (.A(_10831_),
    .B(_10832_),
    .Y(_10833_));
 sky130_fd_sc_hd__nor2_2 _33181_ (.A(_10829_),
    .B(_10833_),
    .Y(_10834_));
 sky130_fd_sc_hd__clkbuf_4 _33182_ (.A(\pcpi_mul.rs2[29] ),
    .X(_10835_));
 sky130_fd_sc_hd__buf_2 _33183_ (.A(_10835_),
    .X(_10836_));
 sky130_fd_sc_hd__a22oi_4 _33184_ (.A1(_10836_),
    .A2(_06020_),
    .B1(_19587_),
    .B2(_05264_),
    .Y(_10837_));
 sky130_fd_sc_hd__nor2_8 _33185_ (.A(_10820_),
    .B(_10821_),
    .Y(_10838_));
 sky130_fd_sc_hd__o21ai_2 _33186_ (.A1(_10837_),
    .A2(_10838_),
    .B1(_10824_),
    .Y(_10839_));
 sky130_fd_sc_hd__nand3_4 _33187_ (.A(_10826_),
    .B(_10834_),
    .C(_10839_),
    .Y(_10840_));
 sky130_fd_sc_hd__o21ai_2 _33188_ (.A1(_10837_),
    .A2(_10838_),
    .B1(_10825_),
    .Y(_10841_));
 sky130_fd_sc_hd__nand3_4 _33189_ (.A(_10822_),
    .B(_10823_),
    .C(_10824_),
    .Y(_10842_));
 sky130_fd_sc_hd__o211ai_4 _33190_ (.A1(_10829_),
    .A2(_10833_),
    .B1(_10841_),
    .C1(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__nand3b_4 _33191_ (.A_N(_10289_),
    .B(_10840_),
    .C(_10843_),
    .Y(_10844_));
 sky130_fd_sc_hd__nand2_2 _33192_ (.A(_10843_),
    .B(_10840_),
    .Y(_10845_));
 sky130_fd_sc_hd__nand2_4 _33193_ (.A(_10845_),
    .B(_10289_),
    .Y(_10846_));
 sky130_fd_sc_hd__a21o_1 _33194_ (.A1(_10279_),
    .A2(_10277_),
    .B1(_10284_),
    .X(_10847_));
 sky130_fd_sc_hd__a22oi_4 _33195_ (.A1(_09722_),
    .A2(_05383_),
    .B1(_09723_),
    .B2(_05380_),
    .Y(_10848_));
 sky130_fd_sc_hd__nand3_4 _33196_ (.A(_09229_),
    .B(_19599_),
    .C(_05208_),
    .Y(_10849_));
 sky130_fd_sc_hd__nor2_4 _33197_ (.A(_05278_),
    .B(_10849_),
    .Y(_10850_));
 sky130_fd_sc_hd__nand2_2 _33198_ (.A(_19602_),
    .B(_05545_),
    .Y(_10851_));
 sky130_fd_sc_hd__o21ai_2 _33199_ (.A1(_10848_),
    .A2(_10850_),
    .B1(_10851_),
    .Y(_10852_));
 sky130_vsdinv _33200_ (.A(_10851_),
    .Y(_10853_));
 sky130_fd_sc_hd__a22o_2 _33201_ (.A1(_10256_),
    .A2(_19917_),
    .B1(_10257_),
    .B2(_05656_),
    .X(_10854_));
 sky130_fd_sc_hd__o211ai_2 _33202_ (.A1(net452),
    .A2(_10849_),
    .B1(_10853_),
    .C1(_10854_),
    .Y(_10855_));
 sky130_fd_sc_hd__nand3_4 _33203_ (.A(_10847_),
    .B(_10852_),
    .C(_10855_),
    .Y(_10856_));
 sky130_fd_sc_hd__o21ai_2 _33204_ (.A1(_10848_),
    .A2(_10850_),
    .B1(_10853_),
    .Y(_10857_));
 sky130_fd_sc_hd__a21oi_2 _33205_ (.A1(_10279_),
    .A2(_10277_),
    .B1(_10284_),
    .Y(_10858_));
 sky130_fd_sc_hd__o211ai_2 _33206_ (.A1(_05551_),
    .A2(_10849_),
    .B1(_10851_),
    .C1(_10854_),
    .Y(_10859_));
 sky130_fd_sc_hd__nand3_4 _33207_ (.A(_10857_),
    .B(_10858_),
    .C(_10859_),
    .Y(_10860_));
 sky130_fd_sc_hd__a21oi_4 _33208_ (.A1(_10258_),
    .A2(_10255_),
    .B1(_10253_),
    .Y(_10861_));
 sky130_vsdinv _33209_ (.A(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__a21oi_2 _33210_ (.A1(_10856_),
    .A2(_10860_),
    .B1(_10862_),
    .Y(_10863_));
 sky130_fd_sc_hd__nand3_2 _33211_ (.A(_10856_),
    .B(_10860_),
    .C(_10862_),
    .Y(_10864_));
 sky130_vsdinv _33212_ (.A(_10864_),
    .Y(_10865_));
 sky130_fd_sc_hd__o2bb2ai_4 _33213_ (.A1_N(_10844_),
    .A2_N(_10846_),
    .B1(_10863_),
    .B2(_10865_),
    .Y(_10866_));
 sky130_fd_sc_hd__nand2_2 _33214_ (.A(_10860_),
    .B(_10862_),
    .Y(_10867_));
 sky130_vsdinv _33215_ (.A(_10856_),
    .Y(_10868_));
 sky130_fd_sc_hd__nand2_1 _33216_ (.A(_10856_),
    .B(_10860_),
    .Y(_10869_));
 sky130_fd_sc_hd__nand2_2 _33217_ (.A(_10869_),
    .B(_10861_),
    .Y(_10870_));
 sky130_fd_sc_hd__o2111ai_4 _33218_ (.A1(_10867_),
    .A2(_10868_),
    .B1(_10870_),
    .C1(_10844_),
    .D1(_10846_),
    .Y(_10871_));
 sky130_fd_sc_hd__a21oi_4 _33219_ (.A1(_10866_),
    .A2(_10871_),
    .B1(_10294_),
    .Y(_10872_));
 sky130_fd_sc_hd__and2_1 _33220_ (.A(_10845_),
    .B(_10289_),
    .X(_10873_));
 sky130_fd_sc_hd__nand3_1 _33221_ (.A(_10844_),
    .B(_10870_),
    .C(_10864_),
    .Y(_10874_));
 sky130_fd_sc_hd__o211a_1 _33222_ (.A1(_10873_),
    .A2(_10874_),
    .B1(_10866_),
    .C1(_10294_),
    .X(_10875_));
 sky130_fd_sc_hd__o2bb2ai_4 _33223_ (.A1_N(_10809_),
    .A2_N(_10819_),
    .B1(_10872_),
    .B2(_10875_),
    .Y(_10876_));
 sky130_fd_sc_hd__nand2_2 _33224_ (.A(_10815_),
    .B(_10818_),
    .Y(_10877_));
 sky130_fd_sc_hd__nand3_4 _33225_ (.A(_10294_),
    .B(_10866_),
    .C(_10871_),
    .Y(_10878_));
 sky130_fd_sc_hd__o2bb2ai_4 _33226_ (.A1_N(_10871_),
    .A2_N(_10866_),
    .B1(_10290_),
    .B2(_10296_),
    .Y(_10879_));
 sky130_fd_sc_hd__o2111ai_4 _33227_ (.A1(_10808_),
    .A2(_10877_),
    .B1(_10878_),
    .C1(_10809_),
    .D1(_10879_),
    .Y(_10880_));
 sky130_fd_sc_hd__nand3_4 _33228_ (.A(_10295_),
    .B(_10336_),
    .C(_10341_),
    .Y(_10881_));
 sky130_fd_sc_hd__nand2_4 _33229_ (.A(_10881_),
    .B(_10299_),
    .Y(_10882_));
 sky130_fd_sc_hd__a21oi_4 _33230_ (.A1(_10876_),
    .A2(_10880_),
    .B1(_10882_),
    .Y(_10883_));
 sky130_fd_sc_hd__nand3_1 _33231_ (.A(_10809_),
    .B(_10819_),
    .C(_10878_),
    .Y(_10884_));
 sky130_fd_sc_hd__o211a_4 _33232_ (.A1(_10872_),
    .A2(_10884_),
    .B1(_10876_),
    .C1(_10882_),
    .X(_10885_));
 sky130_fd_sc_hd__o22ai_4 _33233_ (.A1(_10774_),
    .A2(_10776_),
    .B1(_10883_),
    .B2(_10885_),
    .Y(_10886_));
 sky130_vsdinv _33234_ (.A(_10765_),
    .Y(_10887_));
 sky130_fd_sc_hd__nand2_1 _33235_ (.A(_10771_),
    .B(_10773_),
    .Y(_10888_));
 sky130_fd_sc_hd__o2bb2ai_4 _33236_ (.A1_N(_10771_),
    .A2_N(_10765_),
    .B1(_10414_),
    .B2(_10772_),
    .Y(_10889_));
 sky130_fd_sc_hd__nand3_4 _33237_ (.A(_10882_),
    .B(_10876_),
    .C(_10880_),
    .Y(_10890_));
 sky130_fd_sc_hd__a22oi_4 _33238_ (.A1(_10809_),
    .A2(_10819_),
    .B1(_10879_),
    .B2(_10878_),
    .Y(_10891_));
 sky130_fd_sc_hd__o2111a_1 _33239_ (.A1(_10808_),
    .A2(_10877_),
    .B1(_10878_),
    .C1(_10809_),
    .D1(_10879_),
    .X(_10892_));
 sky130_fd_sc_hd__o31a_1 _33240_ (.A1(_10060_),
    .A2(_10291_),
    .A3(_10294_),
    .B1(_10881_),
    .X(_10893_));
 sky130_fd_sc_hd__o21ai_4 _33241_ (.A1(_10891_),
    .A2(_10892_),
    .B1(_10893_),
    .Y(_10894_));
 sky130_fd_sc_hd__o2111ai_4 _33242_ (.A1(_10887_),
    .A2(_10888_),
    .B1(_10889_),
    .C1(_10890_),
    .D1(_10894_),
    .Y(_10895_));
 sky130_fd_sc_hd__nand3_1 _33243_ (.A(_10412_),
    .B(_10419_),
    .C(_10429_),
    .Y(_10896_));
 sky130_fd_sc_hd__nand3_2 _33244_ (.A(_10441_),
    .B(_10347_),
    .C(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__nand2_2 _33245_ (.A(_10897_),
    .B(_10352_),
    .Y(_10898_));
 sky130_fd_sc_hd__a21oi_4 _33246_ (.A1(_10886_),
    .A2(_10895_),
    .B1(_10898_),
    .Y(_10899_));
 sky130_fd_sc_hd__nand3_4 _33247_ (.A(_10890_),
    .B(_10889_),
    .C(_10775_),
    .Y(_10900_));
 sky130_fd_sc_hd__o211a_2 _33248_ (.A1(_10883_),
    .A2(_10900_),
    .B1(_10886_),
    .C1(_10898_),
    .X(_10901_));
 sky130_fd_sc_hd__o22ai_4 _33249_ (.A1(_10696_),
    .A2(_10699_),
    .B1(_10899_),
    .B2(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__nand3_4 _33250_ (.A(_10898_),
    .B(_10886_),
    .C(_10895_),
    .Y(_10903_));
 sky130_fd_sc_hd__and3_2 _33251_ (.A(_10690_),
    .B(_10691_),
    .C(_10692_),
    .X(_10904_));
 sky130_fd_sc_hd__o22ai_4 _33252_ (.A1(_10485_),
    .A2(_10694_),
    .B1(_10697_),
    .B2(_10904_),
    .Y(_10905_));
 sky130_fd_sc_hd__a22oi_4 _33253_ (.A1(_10889_),
    .A2(_10775_),
    .B1(_10894_),
    .B2(_10890_),
    .Y(_10906_));
 sky130_fd_sc_hd__nor2_2 _33254_ (.A(_10883_),
    .B(_10900_),
    .Y(_10907_));
 sky130_fd_sc_hd__nand2_1 _33255_ (.A(_10349_),
    .B(_10351_),
    .Y(_10908_));
 sky130_fd_sc_hd__o21a_1 _33256_ (.A1(_10908_),
    .A2(_10344_),
    .B1(_10897_),
    .X(_10909_));
 sky130_fd_sc_hd__o21ai_4 _33257_ (.A1(_10906_),
    .A2(_10907_),
    .B1(_10909_),
    .Y(_10910_));
 sky130_fd_sc_hd__o2111ai_4 _33258_ (.A1(_10697_),
    .A2(_10698_),
    .B1(_10903_),
    .C1(_10905_),
    .D1(_10910_),
    .Y(_10911_));
 sky130_fd_sc_hd__a21oi_2 _33259_ (.A1(_10426_),
    .A2(_10431_),
    .B1(_10249_),
    .Y(_10912_));
 sky130_fd_sc_hd__a31oi_4 _33260_ (.A1(_10432_),
    .A2(_10545_),
    .A3(_10547_),
    .B1(_10912_),
    .Y(_10913_));
 sky130_fd_sc_hd__nand3_4 _33261_ (.A(_10902_),
    .B(_10911_),
    .C(_10913_),
    .Y(_10914_));
 sky130_fd_sc_hd__nand2_1 _33262_ (.A(_10688_),
    .B(_10693_),
    .Y(_10915_));
 sky130_fd_sc_hd__nand2_4 _33263_ (.A(_10915_),
    .B(_10695_),
    .Y(_10916_));
 sky130_fd_sc_hd__or2_2 _33264_ (.A(_10485_),
    .B(_10694_),
    .X(_10917_));
 sky130_fd_sc_hd__nand3_4 _33265_ (.A(_10917_),
    .B(_10688_),
    .C(_10693_),
    .Y(_10918_));
 sky130_fd_sc_hd__o2bb2ai_2 _33266_ (.A1_N(_10916_),
    .A2_N(_10918_),
    .B1(_10899_),
    .B2(_10901_),
    .Y(_10919_));
 sky130_fd_sc_hd__nand2_1 _33267_ (.A(_10917_),
    .B(_10688_),
    .Y(_10920_));
 sky130_fd_sc_hd__o2111ai_4 _33268_ (.A1(_10904_),
    .A2(_10920_),
    .B1(_10903_),
    .C1(_10916_),
    .D1(_10910_),
    .Y(_10921_));
 sky130_fd_sc_hd__nand3_1 _33269_ (.A(_10432_),
    .B(_10545_),
    .C(_10547_),
    .Y(_10922_));
 sky130_fd_sc_hd__nand2_1 _33270_ (.A(_10922_),
    .B(_10443_),
    .Y(_10923_));
 sky130_fd_sc_hd__nand3_4 _33271_ (.A(_10919_),
    .B(_10921_),
    .C(_10923_),
    .Y(_10924_));
 sky130_vsdinv _33272_ (.A(_10519_),
    .Y(_10925_));
 sky130_fd_sc_hd__nor2_8 _33273_ (.A(_10523_),
    .B(_10925_),
    .Y(_10926_));
 sky130_vsdinv _33274_ (.A(_10926_),
    .Y(_10927_));
 sky130_fd_sc_hd__and2_2 _33275_ (.A(_10551_),
    .B(_10546_),
    .X(_10928_));
 sky130_fd_sc_hd__nor2_1 _33276_ (.A(_10927_),
    .B(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__nand2_2 _33277_ (.A(_10551_),
    .B(_10546_),
    .Y(_10930_));
 sky130_fd_sc_hd__nor2_1 _33278_ (.A(_10926_),
    .B(_10930_),
    .Y(_10931_));
 sky130_fd_sc_hd__o2bb2ai_2 _33279_ (.A1_N(_10914_),
    .A2_N(_10924_),
    .B1(_10929_),
    .B2(_10931_),
    .Y(_10932_));
 sky130_fd_sc_hd__a21boi_2 _33280_ (.A1(_10561_),
    .A2(_10564_),
    .B1_N(_10553_),
    .Y(_10933_));
 sky130_fd_sc_hd__nor2_4 _33281_ (.A(_10927_),
    .B(_10930_),
    .Y(_10934_));
 sky130_fd_sc_hd__nor2_8 _33282_ (.A(_10926_),
    .B(_10928_),
    .Y(_10935_));
 sky130_fd_sc_hd__nor2_4 _33283_ (.A(_10934_),
    .B(_10935_),
    .Y(_10936_));
 sky130_fd_sc_hd__nand3b_4 _33284_ (.A_N(_10936_),
    .B(_10914_),
    .C(_10924_),
    .Y(_10937_));
 sky130_fd_sc_hd__nand3_4 _33285_ (.A(_10932_),
    .B(_10933_),
    .C(_10937_),
    .Y(_10938_));
 sky130_fd_sc_hd__o2bb2ai_2 _33286_ (.A1_N(_10914_),
    .A2_N(_10924_),
    .B1(_10935_),
    .B2(_10934_),
    .Y(_10939_));
 sky130_vsdinv _33287_ (.A(_10549_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand2_1 _33288_ (.A(_10247_),
    .B(_10552_),
    .Y(_10941_));
 sky130_fd_sc_hd__o2bb2ai_2 _33289_ (.A1_N(_10561_),
    .A2_N(_10564_),
    .B1(_10940_),
    .B2(_10941_),
    .Y(_10942_));
 sky130_fd_sc_hd__nand3_2 _33290_ (.A(_10924_),
    .B(_10914_),
    .C(_10936_),
    .Y(_10943_));
 sky130_fd_sc_hd__nand3_4 _33291_ (.A(_10939_),
    .B(_10942_),
    .C(_10943_),
    .Y(_10944_));
 sky130_fd_sc_hd__nand3_4 _33292_ (.A(_10938_),
    .B(_10944_),
    .C(_10568_),
    .Y(_10945_));
 sky130_fd_sc_hd__nand2_2 _33293_ (.A(_10577_),
    .B(_10224_),
    .Y(_10946_));
 sky130_vsdinv _33294_ (.A(_10568_),
    .Y(_10947_));
 sky130_fd_sc_hd__nand2_1 _33295_ (.A(_10938_),
    .B(_10944_),
    .Y(_10948_));
 sky130_fd_sc_hd__a22oi_4 _33296_ (.A1(_10946_),
    .A2(_10571_),
    .B1(_10947_),
    .B2(_10948_),
    .Y(_10949_));
 sky130_fd_sc_hd__o2bb2ai_4 _33297_ (.A1_N(_10944_),
    .A2_N(_10938_),
    .B1(_10566_),
    .B2(_10567_),
    .Y(_10950_));
 sky130_fd_sc_hd__nand2_2 _33298_ (.A(_10946_),
    .B(_10571_),
    .Y(_10951_));
 sky130_fd_sc_hd__a21oi_4 _33299_ (.A1(_10950_),
    .A2(_10945_),
    .B1(_10951_),
    .Y(_10952_));
 sky130_fd_sc_hd__a21oi_4 _33300_ (.A1(_10945_),
    .A2(_10949_),
    .B1(_10952_),
    .Y(_10953_));
 sky130_fd_sc_hd__nor2_1 _33301_ (.A(_10584_),
    .B(_10592_),
    .Y(_10954_));
 sky130_fd_sc_hd__xnor2_1 _33302_ (.A(_10953_),
    .B(_10954_),
    .Y(_02650_));
 sky130_fd_sc_hd__nand2_4 _33303_ (.A(_10895_),
    .B(_10890_),
    .Y(_10955_));
 sky130_fd_sc_hd__nor2_2 _33304_ (.A(_10727_),
    .B(_10723_),
    .Y(_10956_));
 sky130_fd_sc_hd__buf_6 _33305_ (.A(_08061_),
    .X(_10957_));
 sky130_fd_sc_hd__a22oi_4 _33306_ (.A1(net445),
    .A2(_19874_),
    .B1(_06423_),
    .B2(_10957_),
    .Y(_10958_));
 sky130_vsdinv _33307_ (.A(_07556_),
    .Y(_10959_));
 sky130_fd_sc_hd__buf_8 _33308_ (.A(_10959_),
    .X(_10960_));
 sky130_fd_sc_hd__nand3_4 _33309_ (.A(_06606_),
    .B(_06898_),
    .C(_08735_),
    .Y(_10961_));
 sky130_fd_sc_hd__nor2_8 _33310_ (.A(_10960_),
    .B(_10961_),
    .Y(_10962_));
 sky130_fd_sc_hd__nand2_2 _33311_ (.A(_06419_),
    .B(_07705_),
    .Y(_10963_));
 sky130_fd_sc_hd__o21ai_2 _33312_ (.A1(_10958_),
    .A2(_10962_),
    .B1(_10963_),
    .Y(_10964_));
 sky130_fd_sc_hd__a22o_2 _33313_ (.A1(_06342_),
    .A2(_10733_),
    .B1(_06343_),
    .B2(_10957_),
    .X(_10965_));
 sky130_vsdinv _33314_ (.A(_10963_),
    .Y(_10966_));
 sky130_fd_sc_hd__nand3b_2 _33315_ (.A_N(_10962_),
    .B(_10965_),
    .C(_10966_),
    .Y(_10967_));
 sky130_fd_sc_hd__o211ai_4 _33316_ (.A1(_10726_),
    .A2(_10956_),
    .B1(_10964_),
    .C1(_10967_),
    .Y(_10968_));
 sky130_fd_sc_hd__o21ai_4 _33317_ (.A1(_10958_),
    .A2(_10962_),
    .B1(_10966_),
    .Y(_10969_));
 sky130_fd_sc_hd__a21oi_4 _33318_ (.A1(_10734_),
    .A2(_10728_),
    .B1(_10726_),
    .Y(_10970_));
 sky130_fd_sc_hd__buf_4 _33319_ (.A(_10959_),
    .X(_10971_));
 sky130_fd_sc_hd__o211ai_4 _33320_ (.A1(_10971_),
    .A2(_10961_),
    .B1(_10963_),
    .C1(_10965_),
    .Y(_10972_));
 sky130_fd_sc_hd__nand3_4 _33321_ (.A(_10969_),
    .B(_10970_),
    .C(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__nand2_1 _33322_ (.A(_10968_),
    .B(_10973_),
    .Y(_10974_));
 sky130_fd_sc_hd__a22oi_4 _33323_ (.A1(_06327_),
    .A2(_19866_),
    .B1(_05737_),
    .B2(_19863_),
    .Y(_10975_));
 sky130_fd_sc_hd__nand2_2 _33324_ (.A(_06883_),
    .B(_08056_),
    .Y(_10976_));
 sky130_fd_sc_hd__nand2_1 _33325_ (.A(_06399_),
    .B(_08332_),
    .Y(_10977_));
 sky130_fd_sc_hd__nor2_2 _33326_ (.A(_10976_),
    .B(_10977_),
    .Y(_10978_));
 sky130_fd_sc_hd__nand2_2 _33327_ (.A(_05732_),
    .B(_09082_),
    .Y(_10979_));
 sky130_fd_sc_hd__o21bai_2 _33328_ (.A1(_10975_),
    .A2(_10978_),
    .B1_N(_10979_),
    .Y(_10980_));
 sky130_fd_sc_hd__buf_4 _33329_ (.A(_10458_),
    .X(_10981_));
 sky130_fd_sc_hd__nand3b_4 _33330_ (.A_N(_10976_),
    .B(_06160_),
    .C(_10981_),
    .Y(_10982_));
 sky130_fd_sc_hd__nand2_2 _33331_ (.A(_10976_),
    .B(_10977_),
    .Y(_10983_));
 sky130_fd_sc_hd__nand3_4 _33332_ (.A(_10982_),
    .B(_10979_),
    .C(_10983_),
    .Y(_10984_));
 sky130_fd_sc_hd__nand2_4 _33333_ (.A(_10980_),
    .B(_10984_),
    .Y(_10985_));
 sky130_fd_sc_hd__and2_1 _33334_ (.A(_10974_),
    .B(_10985_),
    .X(_10986_));
 sky130_fd_sc_hd__nor2_2 _33335_ (.A(_10985_),
    .B(_10974_),
    .Y(_10987_));
 sky130_fd_sc_hd__nand2_2 _33336_ (.A(_10796_),
    .B(_10797_),
    .Y(_10988_));
 sky130_fd_sc_hd__a21oi_4 _33337_ (.A1(_10800_),
    .A2(_10988_),
    .B1(_10798_),
    .Y(_10989_));
 sky130_fd_sc_hd__buf_6 _33338_ (.A(_06924_),
    .X(_10990_));
 sky130_fd_sc_hd__buf_6 _33339_ (.A(_08623_),
    .X(_10991_));
 sky130_fd_sc_hd__a22oi_4 _33340_ (.A1(_10990_),
    .A2(_07060_),
    .B1(_10991_),
    .B2(_06804_),
    .Y(_10992_));
 sky130_fd_sc_hd__clkinv_8 _33341_ (.A(_06803_),
    .Y(_10993_));
 sky130_fd_sc_hd__nor2_4 _33342_ (.A(_10993_),
    .B(_10700_),
    .Y(_10994_));
 sky130_fd_sc_hd__nand2_2 _33343_ (.A(_07435_),
    .B(_08734_),
    .Y(_10995_));
 sky130_vsdinv _33344_ (.A(_10995_),
    .Y(_10996_));
 sky130_fd_sc_hd__o21ai_2 _33345_ (.A1(_10992_),
    .A2(_10994_),
    .B1(_10996_),
    .Y(_10997_));
 sky130_fd_sc_hd__buf_4 _33346_ (.A(_08190_),
    .X(_10998_));
 sky130_fd_sc_hd__clkbuf_4 _33347_ (.A(_07928_),
    .X(_10999_));
 sky130_fd_sc_hd__a22o_2 _33348_ (.A1(_10998_),
    .A2(_06635_),
    .B1(_10999_),
    .B2(_07055_),
    .X(_11000_));
 sky130_fd_sc_hd__o211ai_4 _33349_ (.A1(_10993_),
    .A2(_10700_),
    .B1(_10995_),
    .C1(_11000_),
    .Y(_11001_));
 sky130_fd_sc_hd__nand3_4 _33350_ (.A(_10989_),
    .B(_10997_),
    .C(_11001_),
    .Y(_11002_));
 sky130_fd_sc_hd__buf_4 _33351_ (.A(_10364_),
    .X(_11003_));
 sky130_fd_sc_hd__a31o_1 _33352_ (.A1(_10988_),
    .A2(_11003_),
    .A3(_19892_),
    .B1(_10798_),
    .X(_11004_));
 sky130_fd_sc_hd__nand3b_2 _33353_ (.A_N(_10994_),
    .B(_11000_),
    .C(_10996_),
    .Y(_11005_));
 sky130_fd_sc_hd__o21ai_2 _33354_ (.A1(_10992_),
    .A2(_10994_),
    .B1(_10995_),
    .Y(_11006_));
 sky130_fd_sc_hd__nand3_4 _33355_ (.A(_11004_),
    .B(_11005_),
    .C(_11006_),
    .Y(_11007_));
 sky130_vsdinv _33356_ (.A(_10701_),
    .Y(_11008_));
 sky130_fd_sc_hd__nor2_2 _33357_ (.A(_10704_),
    .B(_10706_),
    .Y(_11009_));
 sky130_fd_sc_hd__o2bb2ai_4 _33358_ (.A1_N(_11002_),
    .A2_N(_11007_),
    .B1(_11008_),
    .B2(_11009_),
    .Y(_11010_));
 sky130_fd_sc_hd__and3_1 _33359_ (.A(_10701_),
    .B(net458),
    .C(_19882_),
    .X(_11011_));
 sky130_fd_sc_hd__o211ai_4 _33360_ (.A1(_10706_),
    .A2(_11011_),
    .B1(_11002_),
    .C1(_11007_),
    .Y(_11012_));
 sky130_fd_sc_hd__nand2_1 _33361_ (.A(_10709_),
    .B(_10716_),
    .Y(_11013_));
 sky130_fd_sc_hd__nand2_4 _33362_ (.A(_11013_),
    .B(_10712_),
    .Y(_11014_));
 sky130_fd_sc_hd__a21oi_4 _33363_ (.A1(_11010_),
    .A2(_11012_),
    .B1(_11014_),
    .Y(_11015_));
 sky130_fd_sc_hd__a21oi_2 _33364_ (.A1(_10705_),
    .A2(_10707_),
    .B1(_10708_),
    .Y(_11016_));
 sky130_fd_sc_hd__o211a_4 _33365_ (.A1(_11016_),
    .A2(_10720_),
    .B1(_11012_),
    .C1(_11010_),
    .X(_11017_));
 sky130_fd_sc_hd__o22ai_4 _33366_ (.A1(_10986_),
    .A2(_10987_),
    .B1(_11015_),
    .B2(_11017_),
    .Y(_11018_));
 sky130_fd_sc_hd__a21o_1 _33367_ (.A1(_11010_),
    .A2(_11012_),
    .B1(_11014_),
    .X(_11019_));
 sky130_fd_sc_hd__nand3_4 _33368_ (.A(_11014_),
    .B(_11010_),
    .C(_11012_),
    .Y(_11020_));
 sky130_fd_sc_hd__a21oi_4 _33369_ (.A1(_10969_),
    .A2(_10972_),
    .B1(_10970_),
    .Y(_11021_));
 sky130_fd_sc_hd__nand2_2 _33370_ (.A(_10973_),
    .B(_10985_),
    .Y(_11022_));
 sky130_fd_sc_hd__a21o_1 _33371_ (.A1(_10968_),
    .A2(_10973_),
    .B1(_10985_),
    .X(_11023_));
 sky130_fd_sc_hd__o21ai_4 _33372_ (.A1(_11021_),
    .A2(_11022_),
    .B1(_11023_),
    .Y(_11024_));
 sky130_fd_sc_hd__nand3_4 _33373_ (.A(_11019_),
    .B(_11020_),
    .C(_11024_),
    .Y(_11025_));
 sky130_fd_sc_hd__a21oi_4 _33374_ (.A1(_10815_),
    .A2(_10818_),
    .B1(_10808_),
    .Y(_11026_));
 sky130_fd_sc_hd__a21oi_4 _33375_ (.A1(_11018_),
    .A2(_11025_),
    .B1(_11026_),
    .Y(_11027_));
 sky130_fd_sc_hd__nand3_4 _33376_ (.A(_11018_),
    .B(_11026_),
    .C(_11025_),
    .Y(_11028_));
 sky130_fd_sc_hd__o21ai_4 _33377_ (.A1(_10756_),
    .A2(_10719_),
    .B1(_10760_),
    .Y(_11029_));
 sky130_fd_sc_hd__nand2_2 _33378_ (.A(_11028_),
    .B(_11029_),
    .Y(_11030_));
 sky130_fd_sc_hd__nor2_2 _33379_ (.A(_11027_),
    .B(_11030_),
    .Y(_11031_));
 sky130_fd_sc_hd__o21a_1 _33380_ (.A1(_11021_),
    .A2(_11022_),
    .B1(_11023_),
    .X(_11032_));
 sky130_fd_sc_hd__nand2_1 _33381_ (.A(_11032_),
    .B(_11020_),
    .Y(_11033_));
 sky130_vsdinv _33382_ (.A(_10818_),
    .Y(_11034_));
 sky130_fd_sc_hd__o21ai_2 _33383_ (.A1(_11034_),
    .A2(_10807_),
    .B1(_10816_),
    .Y(_11035_));
 sky130_fd_sc_hd__o21ai_2 _33384_ (.A1(_11015_),
    .A2(_11017_),
    .B1(_11024_),
    .Y(_11036_));
 sky130_fd_sc_hd__o211ai_4 _33385_ (.A1(_11015_),
    .A2(_11033_),
    .B1(_11035_),
    .C1(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__a21oi_4 _33386_ (.A1(_11037_),
    .A2(_11028_),
    .B1(_11029_),
    .Y(_11038_));
 sky130_fd_sc_hd__a31o_1 _33387_ (.A1(_10783_),
    .A2(_19617_),
    .A3(_19902_),
    .B1(_10781_),
    .X(_11039_));
 sky130_fd_sc_hd__nand2_4 _33388_ (.A(_19615_),
    .B(_05976_),
    .Y(_11040_));
 sky130_vsdinv _33389_ (.A(_11040_),
    .Y(_11041_));
 sky130_fd_sc_hd__a22o_1 _33390_ (.A1(_10073_),
    .A2(_06264_),
    .B1(_09680_),
    .B2(_07789_),
    .X(_11042_));
 sky130_fd_sc_hd__o211ai_2 _33391_ (.A1(_06272_),
    .A2(_10791_),
    .B1(_11041_),
    .C1(_11042_),
    .Y(_11043_));
 sky130_fd_sc_hd__a22oi_4 _33392_ (.A1(_10073_),
    .A2(_05673_),
    .B1(_10066_),
    .B2(_06441_),
    .Y(_11044_));
 sky130_fd_sc_hd__nor2_4 _33393_ (.A(net446),
    .B(_10791_),
    .Y(_11045_));
 sky130_fd_sc_hd__o21ai_2 _33394_ (.A1(_11044_),
    .A2(_11045_),
    .B1(_11040_),
    .Y(_11046_));
 sky130_fd_sc_hd__nand3_4 _33395_ (.A(_11039_),
    .B(_11043_),
    .C(_11046_),
    .Y(_11047_));
 sky130_fd_sc_hd__o21ai_2 _33396_ (.A1(_11044_),
    .A2(_11045_),
    .B1(_11041_),
    .Y(_11048_));
 sky130_fd_sc_hd__o21ai_2 _33397_ (.A1(_10787_),
    .A2(_10781_),
    .B1(_10783_),
    .Y(_11049_));
 sky130_fd_sc_hd__o211ai_2 _33398_ (.A1(_06272_),
    .A2(_10791_),
    .B1(_11040_),
    .C1(_11042_),
    .Y(_11050_));
 sky130_fd_sc_hd__nand3_4 _33399_ (.A(_11048_),
    .B(_11049_),
    .C(_11050_),
    .Y(_11051_));
 sky130_fd_sc_hd__nand2_1 _33400_ (.A(_11047_),
    .B(_11051_),
    .Y(_11052_));
 sky130_fd_sc_hd__nand2_1 _33401_ (.A(_10364_),
    .B(_07064_),
    .Y(_11053_));
 sky130_vsdinv _33402_ (.A(_11053_),
    .Y(_11054_));
 sky130_fd_sc_hd__a22oi_4 _33403_ (.A1(_19622_),
    .A2(_06289_),
    .B1(_08565_),
    .B2(_06286_),
    .Y(_11055_));
 sky130_fd_sc_hd__nand2_2 _33404_ (.A(_07757_),
    .B(_05962_),
    .Y(_11056_));
 sky130_fd_sc_hd__nand2_4 _33405_ (.A(_08567_),
    .B(_07281_),
    .Y(_11057_));
 sky130_fd_sc_hd__nor2_8 _33406_ (.A(_11056_),
    .B(_11057_),
    .Y(_11058_));
 sky130_fd_sc_hd__nor3_1 _33407_ (.A(_11054_),
    .B(_11055_),
    .C(_11058_),
    .Y(_11059_));
 sky130_fd_sc_hd__o21ai_2 _33408_ (.A1(_11055_),
    .A2(_11058_),
    .B1(_11054_),
    .Y(_11060_));
 sky130_fd_sc_hd__and2b_2 _33409_ (.A_N(_11059_),
    .B(_11060_),
    .X(_11061_));
 sky130_fd_sc_hd__nand2_4 _33410_ (.A(_11052_),
    .B(_11061_),
    .Y(_11062_));
 sky130_fd_sc_hd__nor2_1 _33411_ (.A(_11055_),
    .B(_11058_),
    .Y(_11063_));
 sky130_fd_sc_hd__nand2_1 _33412_ (.A(_11063_),
    .B(_11053_),
    .Y(_11064_));
 sky130_fd_sc_hd__nand2_4 _33413_ (.A(_11064_),
    .B(_11060_),
    .Y(_11065_));
 sky130_fd_sc_hd__nand3_4 _33414_ (.A(_11065_),
    .B(_11047_),
    .C(_11051_),
    .Y(_11066_));
 sky130_fd_sc_hd__nand2_4 _33415_ (.A(_10867_),
    .B(_10856_),
    .Y(_11067_));
 sky130_fd_sc_hd__a21o_2 _33416_ (.A1(_11062_),
    .A2(_11066_),
    .B1(_11067_),
    .X(_11068_));
 sky130_fd_sc_hd__nand3_4 _33417_ (.A(_11062_),
    .B(_11067_),
    .C(_11066_),
    .Y(_11069_));
 sky130_fd_sc_hd__nand2_1 _33418_ (.A(_10802_),
    .B(_10789_),
    .Y(_11070_));
 sky130_fd_sc_hd__nand2_2 _33419_ (.A(_11070_),
    .B(_10804_),
    .Y(_11071_));
 sky130_fd_sc_hd__a21oi_2 _33420_ (.A1(_11068_),
    .A2(_11069_),
    .B1(_11071_),
    .Y(_11072_));
 sky130_fd_sc_hd__nand3_2 _33421_ (.A(_11068_),
    .B(_11069_),
    .C(_11071_),
    .Y(_11073_));
 sky130_vsdinv _33422_ (.A(_11073_),
    .Y(_11074_));
 sky130_fd_sc_hd__buf_6 _33423_ (.A(\pcpi_mul.rs2[32] ),
    .X(_11075_));
 sky130_fd_sc_hd__nand3_4 _33424_ (.A(_11075_),
    .B(_19575_),
    .C(_19929_),
    .Y(_11076_));
 sky130_fd_sc_hd__nor2_4 _33425_ (.A(_05198_),
    .B(_11076_),
    .Y(_11077_));
 sky130_fd_sc_hd__buf_4 _33426_ (.A(\pcpi_mul.rs2[31] ),
    .X(_11078_));
 sky130_fd_sc_hd__buf_6 _33427_ (.A(_11078_),
    .X(_11079_));
 sky130_fd_sc_hd__buf_6 _33428_ (.A(_11075_),
    .X(_11080_));
 sky130_fd_sc_hd__a22oi_4 _33429_ (.A1(_11079_),
    .A2(_19930_),
    .B1(_04840_),
    .B2(_11080_),
    .Y(_11081_));
 sky130_fd_sc_hd__nand2_4 _33430_ (.A(_10827_),
    .B(_07828_),
    .Y(_11082_));
 sky130_vsdinv _33431_ (.A(_11082_),
    .Y(_11083_));
 sky130_fd_sc_hd__o21ai_2 _33432_ (.A1(_11077_),
    .A2(_11081_),
    .B1(_11083_),
    .Y(_11084_));
 sky130_vsdinv _33433_ (.A(_10833_),
    .Y(_11085_));
 sky130_fd_sc_hd__nand2_1 _33434_ (.A(_10830_),
    .B(_05441_),
    .Y(_11086_));
 sky130_fd_sc_hd__o21ai_4 _33435_ (.A1(_05198_),
    .A2(_18474_),
    .B1(_11086_),
    .Y(_11087_));
 sky130_fd_sc_hd__o211ai_4 _33436_ (.A1(_05406_),
    .A2(_11076_),
    .B1(_11082_),
    .C1(_11087_),
    .Y(_11088_));
 sky130_fd_sc_hd__nand3_4 _33437_ (.A(_11084_),
    .B(_11085_),
    .C(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__nand3b_2 _33438_ (.A_N(_11077_),
    .B(_11083_),
    .C(_11087_),
    .Y(_11090_));
 sky130_fd_sc_hd__nand2_2 _33439_ (.A(_11090_),
    .B(_10833_),
    .Y(_11091_));
 sky130_fd_sc_hd__nand2_1 _33440_ (.A(_11089_),
    .B(_11091_),
    .Y(_11092_));
 sky130_fd_sc_hd__a22oi_4 _33441_ (.A1(_19583_),
    .A2(_05838_),
    .B1(_10282_),
    .B2(_06330_),
    .Y(_11093_));
 sky130_fd_sc_hd__buf_2 _33442_ (.A(\pcpi_mul.rs2[28] ),
    .X(_11094_));
 sky130_fd_sc_hd__nand3_4 _33443_ (.A(net469),
    .B(net494),
    .C(_19920_),
    .Y(_11095_));
 sky130_fd_sc_hd__nor2_2 _33444_ (.A(_05154_),
    .B(_11095_),
    .Y(_11096_));
 sky130_fd_sc_hd__nand2_2 _33445_ (.A(_10251_),
    .B(_05378_),
    .Y(_11097_));
 sky130_vsdinv _33446_ (.A(_11097_),
    .Y(_11098_));
 sky130_fd_sc_hd__o21ai_2 _33447_ (.A1(_11093_),
    .A2(_11096_),
    .B1(_11098_),
    .Y(_11099_));
 sky130_fd_sc_hd__a22o_2 _33448_ (.A1(_10281_),
    .A2(_19924_),
    .B1(_10282_),
    .B2(_06330_),
    .X(_11100_));
 sky130_fd_sc_hd__o211ai_4 _33449_ (.A1(_05155_),
    .A2(_11095_),
    .B1(_11097_),
    .C1(_11100_),
    .Y(_11101_));
 sky130_fd_sc_hd__and2_1 _33450_ (.A(_11099_),
    .B(_11101_),
    .X(_11102_));
 sky130_fd_sc_hd__nand2_1 _33451_ (.A(_11092_),
    .B(_11102_),
    .Y(_11103_));
 sky130_vsdinv _33452_ (.A(_10840_),
    .Y(_11104_));
 sky130_fd_sc_hd__nand2_4 _33453_ (.A(_11099_),
    .B(_11101_),
    .Y(_11105_));
 sky130_fd_sc_hd__nand3_4 _33454_ (.A(_11089_),
    .B(_11091_),
    .C(_11105_),
    .Y(_11106_));
 sky130_fd_sc_hd__nand3_4 _33455_ (.A(_11103_),
    .B(_11104_),
    .C(_11106_),
    .Y(_11107_));
 sky130_fd_sc_hd__nand2_1 _33456_ (.A(_11092_),
    .B(_11105_),
    .Y(_11108_));
 sky130_fd_sc_hd__nand3_2 _33457_ (.A(_11102_),
    .B(_11091_),
    .C(_11089_),
    .Y(_11109_));
 sky130_fd_sc_hd__nand3_4 _33458_ (.A(_11108_),
    .B(_10840_),
    .C(_11109_),
    .Y(_11110_));
 sky130_fd_sc_hd__or2_2 _33459_ (.A(_10853_),
    .B(_10850_),
    .X(_11111_));
 sky130_fd_sc_hd__nand2_4 _33460_ (.A(_09227_),
    .B(_05769_),
    .Y(_11112_));
 sky130_fd_sc_hd__nand3_2 _33461_ (.A(_11112_),
    .B(_10260_),
    .C(_05484_),
    .Y(_11113_));
 sky130_fd_sc_hd__nand2_4 _33462_ (.A(_09229_),
    .B(_19913_),
    .Y(_11114_));
 sky130_fd_sc_hd__nand3_2 _33463_ (.A(_11114_),
    .B(_10261_),
    .C(_05770_),
    .Y(_11115_));
 sky130_fd_sc_hd__o211ai_4 _33464_ (.A1(_08578_),
    .A2(net449),
    .B1(_11113_),
    .C1(_11115_),
    .Y(_11116_));
 sky130_fd_sc_hd__nand3_2 _33465_ (.A(_09722_),
    .B(_10257_),
    .C(_05656_),
    .Y(_11117_));
 sky130_fd_sc_hd__nand2_1 _33466_ (.A(_11114_),
    .B(_11112_),
    .Y(_11118_));
 sky130_fd_sc_hd__o2111ai_4 _33467_ (.A1(_08197_),
    .A2(_11117_),
    .B1(_19603_),
    .C1(_06106_),
    .D1(_11118_),
    .Y(_11119_));
 sky130_fd_sc_hd__nor2_1 _33468_ (.A(_10825_),
    .B(_10838_),
    .Y(_11120_));
 sky130_fd_sc_hd__o2bb2ai_1 _33469_ (.A1_N(_11116_),
    .A2_N(_11119_),
    .B1(_10837_),
    .B2(_11120_),
    .Y(_11121_));
 sky130_fd_sc_hd__a21oi_2 _33470_ (.A1(_10820_),
    .A2(_10821_),
    .B1(_10824_),
    .Y(_11122_));
 sky130_fd_sc_hd__o211ai_4 _33471_ (.A1(_10838_),
    .A2(_11122_),
    .B1(_11116_),
    .C1(_11119_),
    .Y(_11123_));
 sky130_fd_sc_hd__a22oi_4 _33472_ (.A1(_10854_),
    .A2(_11111_),
    .B1(_11121_),
    .B2(_11123_),
    .Y(_11124_));
 sky130_fd_sc_hd__o21ai_2 _33473_ (.A1(_10853_),
    .A2(_10850_),
    .B1(_10854_),
    .Y(_11125_));
 sky130_fd_sc_hd__o21ai_2 _33474_ (.A1(_10820_),
    .A2(_10821_),
    .B1(_10824_),
    .Y(_11126_));
 sky130_fd_sc_hd__a22oi_4 _33475_ (.A1(_10823_),
    .A2(_11126_),
    .B1(_11119_),
    .B2(_11116_),
    .Y(_11127_));
 sky130_fd_sc_hd__nor2_2 _33476_ (.A(_11125_),
    .B(_11127_),
    .Y(_11128_));
 sky130_fd_sc_hd__and2_1 _33477_ (.A(_11128_),
    .B(_11123_),
    .X(_11129_));
 sky130_fd_sc_hd__o2bb2ai_4 _33478_ (.A1_N(_11107_),
    .A2_N(_11110_),
    .B1(_11124_),
    .B2(_11129_),
    .Y(_11130_));
 sky130_fd_sc_hd__a21oi_4 _33479_ (.A1(_11123_),
    .A2(_11128_),
    .B1(_11124_),
    .Y(_11131_));
 sky130_fd_sc_hd__nand3_4 _33480_ (.A(_11107_),
    .B(_11110_),
    .C(_11131_),
    .Y(_11132_));
 sky130_fd_sc_hd__nor2_1 _33481_ (.A(_10289_),
    .B(_10845_),
    .Y(_11133_));
 sky130_fd_sc_hd__a31o_2 _33482_ (.A1(_10846_),
    .A2(_10870_),
    .A3(_10864_),
    .B1(_11133_),
    .X(_11134_));
 sky130_fd_sc_hd__a21oi_4 _33483_ (.A1(_11130_),
    .A2(_11132_),
    .B1(_11134_),
    .Y(_11135_));
 sky130_fd_sc_hd__and3_1 _33484_ (.A(_10846_),
    .B(_10870_),
    .C(_10864_),
    .X(_11136_));
 sky130_fd_sc_hd__o211a_2 _33485_ (.A1(_11133_),
    .A2(_11136_),
    .B1(_11132_),
    .C1(_11130_),
    .X(_11137_));
 sky130_fd_sc_hd__o22ai_4 _33486_ (.A1(_11072_),
    .A2(_11074_),
    .B1(_11135_),
    .B2(_11137_),
    .Y(_11138_));
 sky130_fd_sc_hd__a21oi_2 _33487_ (.A1(_11107_),
    .A2(_11110_),
    .B1(_11131_),
    .Y(_11139_));
 sky130_vsdinv _33488_ (.A(_11106_),
    .Y(_11140_));
 sky130_fd_sc_hd__nand2_1 _33489_ (.A(_11084_),
    .B(_11088_),
    .Y(_11141_));
 sky130_vsdinv _33490_ (.A(_10829_),
    .Y(_11142_));
 sky130_fd_sc_hd__nand2_1 _33491_ (.A(_10842_),
    .B(_10841_),
    .Y(_11143_));
 sky130_fd_sc_hd__o2111ai_4 _33492_ (.A1(_11105_),
    .A2(_11141_),
    .B1(_11142_),
    .C1(_11085_),
    .D1(_11143_),
    .Y(_11144_));
 sky130_fd_sc_hd__o211a_2 _33493_ (.A1(_11140_),
    .A2(_11144_),
    .B1(_11131_),
    .C1(_11110_),
    .X(_11145_));
 sky130_fd_sc_hd__o21bai_4 _33494_ (.A1(_11139_),
    .A2(_11145_),
    .B1_N(_11134_),
    .Y(_11146_));
 sky130_fd_sc_hd__a21oi_4 _33495_ (.A1(_11062_),
    .A2(_11066_),
    .B1(_11067_),
    .Y(_11147_));
 sky130_fd_sc_hd__nand2_1 _33496_ (.A(_11065_),
    .B(_11051_),
    .Y(_11148_));
 sky130_vsdinv _33497_ (.A(_11047_),
    .Y(_11149_));
 sky130_fd_sc_hd__o211a_1 _33498_ (.A1(_11148_),
    .A2(_11149_),
    .B1(_11067_),
    .C1(_11062_),
    .X(_11150_));
 sky130_fd_sc_hd__o21ai_2 _33499_ (.A1(_11147_),
    .A2(_11150_),
    .B1(_11071_),
    .Y(_11151_));
 sky130_fd_sc_hd__and2_1 _33500_ (.A(_11070_),
    .B(_10804_),
    .X(_11152_));
 sky130_fd_sc_hd__nand3_2 _33501_ (.A(_11068_),
    .B(_11069_),
    .C(_11152_),
    .Y(_11153_));
 sky130_fd_sc_hd__nand2_4 _33502_ (.A(_11151_),
    .B(_11153_),
    .Y(_11154_));
 sky130_fd_sc_hd__nand3_4 _33503_ (.A(_11130_),
    .B(_11134_),
    .C(_11132_),
    .Y(_11155_));
 sky130_fd_sc_hd__nand3_4 _33504_ (.A(_11146_),
    .B(_11154_),
    .C(_11155_),
    .Y(_11156_));
 sky130_fd_sc_hd__nand2_4 _33505_ (.A(_10880_),
    .B(_10878_),
    .Y(_11157_));
 sky130_fd_sc_hd__a21oi_4 _33506_ (.A1(_11138_),
    .A2(_11156_),
    .B1(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__o211a_1 _33507_ (.A1(_10875_),
    .A2(_10892_),
    .B1(_11156_),
    .C1(_11138_),
    .X(_11159_));
 sky130_fd_sc_hd__o22ai_4 _33508_ (.A1(_11031_),
    .A2(_11038_),
    .B1(_11158_),
    .B2(_11159_),
    .Y(_11160_));
 sky130_fd_sc_hd__a21oi_2 _33509_ (.A1(_11146_),
    .A2(_11155_),
    .B1(_11154_),
    .Y(_11161_));
 sky130_fd_sc_hd__nand2_2 _33510_ (.A(_11130_),
    .B(_11134_),
    .Y(_11162_));
 sky130_fd_sc_hd__o211a_1 _33511_ (.A1(_11145_),
    .A2(_11162_),
    .B1(_11154_),
    .C1(_11146_),
    .X(_11163_));
 sky130_fd_sc_hd__o21bai_4 _33512_ (.A1(_11161_),
    .A2(_11163_),
    .B1_N(_11157_),
    .Y(_11164_));
 sky130_fd_sc_hd__nand3_4 _33513_ (.A(_11138_),
    .B(_11157_),
    .C(_11156_),
    .Y(_11165_));
 sky130_fd_sc_hd__a21oi_4 _33514_ (.A1(_10759_),
    .A2(_10763_),
    .B1(_10722_),
    .Y(_11166_));
 sky130_fd_sc_hd__a31oi_4 _33515_ (.A1(_11018_),
    .A2(_11026_),
    .A3(_11025_),
    .B1(_11166_),
    .Y(_11167_));
 sky130_fd_sc_hd__a21oi_4 _33516_ (.A1(_11037_),
    .A2(_11167_),
    .B1(_11038_),
    .Y(_11168_));
 sky130_fd_sc_hd__nand3_4 _33517_ (.A(_11164_),
    .B(_11165_),
    .C(_11168_),
    .Y(_11169_));
 sky130_fd_sc_hd__nand3_4 _33518_ (.A(_10955_),
    .B(_11160_),
    .C(_11169_),
    .Y(_11170_));
 sky130_fd_sc_hd__o21ai_2 _33519_ (.A1(_11158_),
    .A2(_11159_),
    .B1(_11168_),
    .Y(_11171_));
 sky130_fd_sc_hd__a31oi_4 _33520_ (.A1(_10894_),
    .A2(_10889_),
    .A3(_10775_),
    .B1(_10885_),
    .Y(_11172_));
 sky130_fd_sc_hd__a21o_1 _33521_ (.A1(_11037_),
    .A2(_11028_),
    .B1(_11029_),
    .X(_11173_));
 sky130_fd_sc_hd__o21ai_4 _33522_ (.A1(_11027_),
    .A2(_11030_),
    .B1(_11173_),
    .Y(_11174_));
 sky130_fd_sc_hd__nand3_2 _33523_ (.A(_11164_),
    .B(_11165_),
    .C(_11174_),
    .Y(_11175_));
 sky130_fd_sc_hd__nand3_4 _33524_ (.A(_11171_),
    .B(_11172_),
    .C(_11175_),
    .Y(_11176_));
 sky130_fd_sc_hd__nand2_2 _33525_ (.A(_11170_),
    .B(_11176_),
    .Y(_11177_));
 sky130_fd_sc_hd__buf_6 _33526_ (.A(_09947_),
    .X(_11178_));
 sky130_fd_sc_hd__buf_6 _33527_ (.A(_19838_),
    .X(_11179_));
 sky130_fd_sc_hd__a22oi_4 _33528_ (.A1(_05791_),
    .A2(_11178_),
    .B1(_05780_),
    .B2(_11179_),
    .Y(_11180_));
 sky130_fd_sc_hd__nand2_4 _33529_ (.A(_05772_),
    .B(_19843_),
    .Y(_11181_));
 sky130_fd_sc_hd__nand2_2 _33530_ (.A(_06659_),
    .B(_09946_),
    .Y(_11182_));
 sky130_fd_sc_hd__nor2_4 _33531_ (.A(_11181_),
    .B(_11182_),
    .Y(_11183_));
 sky130_fd_sc_hd__buf_6 _33532_ (.A(\pcpi_mul.rs1[32] ),
    .X(_11184_));
 sky130_fd_sc_hd__nand2_2 _33533_ (.A(_11184_),
    .B(net495),
    .Y(_11185_));
 sky130_fd_sc_hd__clkbuf_4 _33534_ (.A(_11185_),
    .X(_11186_));
 sky130_fd_sc_hd__o21ai_4 _33535_ (.A1(_11180_),
    .A2(_11183_),
    .B1(_11186_),
    .Y(_11187_));
 sky130_fd_sc_hd__nand3b_4 _33536_ (.A_N(_11181_),
    .B(_19674_),
    .C(_11179_),
    .Y(_11188_));
 sky130_vsdinv _33537_ (.A(_11185_),
    .Y(_11189_));
 sky130_fd_sc_hd__nand2_2 _33538_ (.A(_11181_),
    .B(_11182_),
    .Y(_11190_));
 sky130_fd_sc_hd__nand3_4 _33539_ (.A(_11188_),
    .B(_11189_),
    .C(_11190_),
    .Y(_11191_));
 sky130_fd_sc_hd__nand2_1 _33540_ (.A(_11187_),
    .B(_11191_),
    .Y(_11192_));
 sky130_fd_sc_hd__nor2_2 _33541_ (.A(_10609_),
    .B(_10610_),
    .Y(_11193_));
 sky130_fd_sc_hd__a21oi_4 _33542_ (.A1(_10615_),
    .A2(_10612_),
    .B1(_11193_),
    .Y(_11194_));
 sky130_fd_sc_hd__nand2_2 _33543_ (.A(_11192_),
    .B(_11194_),
    .Y(_11195_));
 sky130_fd_sc_hd__a21o_2 _33544_ (.A1(_10615_),
    .A2(_10612_),
    .B1(_11193_),
    .X(_11196_));
 sky130_fd_sc_hd__nand3_4 _33545_ (.A(_11196_),
    .B(_11187_),
    .C(_11191_),
    .Y(_11197_));
 sky130_fd_sc_hd__nand2_1 _33546_ (.A(_11195_),
    .B(_11197_),
    .Y(_11198_));
 sky130_fd_sc_hd__buf_6 _33547_ (.A(_19829_),
    .X(_11199_));
 sky130_fd_sc_hd__buf_4 _33548_ (.A(_10613_),
    .X(_11200_));
 sky130_fd_sc_hd__a22oi_2 _33549_ (.A1(_19680_),
    .A2(_11199_),
    .B1(_05164_),
    .B2(_11200_),
    .Y(_11201_));
 sky130_fd_sc_hd__buf_4 _33550_ (.A(\pcpi_mul.rs1[30] ),
    .X(_11202_));
 sky130_fd_sc_hd__and4_1 _33551_ (.A(_06281_),
    .B(_05223_),
    .C(_19825_),
    .D(_11202_),
    .X(_11203_));
 sky130_fd_sc_hd__nor2_1 _33552_ (.A(_11201_),
    .B(_11203_),
    .Y(_11204_));
 sky130_vsdinv _33553_ (.A(\pcpi_mul.rs1[29] ),
    .Y(_11205_));
 sky130_fd_sc_hd__clkbuf_8 _33554_ (.A(_11205_),
    .X(_11206_));
 sky130_fd_sc_hd__nor2_1 _33555_ (.A(_05491_),
    .B(_11206_),
    .Y(_11207_));
 sky130_fd_sc_hd__nand2_1 _33556_ (.A(_11204_),
    .B(_11207_),
    .Y(_11208_));
 sky130_fd_sc_hd__o21bai_1 _33557_ (.A1(_11201_),
    .A2(_11203_),
    .B1_N(_11207_),
    .Y(_11209_));
 sky130_fd_sc_hd__and2_1 _33558_ (.A(_11208_),
    .B(_11209_),
    .X(_11210_));
 sky130_fd_sc_hd__nand2_1 _33559_ (.A(_11198_),
    .B(_11210_),
    .Y(_11211_));
 sky130_fd_sc_hd__a21boi_4 _33560_ (.A1(_10607_),
    .A2(_10624_),
    .B1_N(_10621_),
    .Y(_11212_));
 sky130_fd_sc_hd__nand2_2 _33561_ (.A(_11208_),
    .B(_11209_),
    .Y(_11213_));
 sky130_fd_sc_hd__nand3_2 _33562_ (.A(_11195_),
    .B(_11197_),
    .C(_11213_),
    .Y(_11214_));
 sky130_fd_sc_hd__nand3_4 _33563_ (.A(_11211_),
    .B(_11212_),
    .C(_11214_),
    .Y(_11215_));
 sky130_fd_sc_hd__nand2_1 _33564_ (.A(_11198_),
    .B(_11213_),
    .Y(_11216_));
 sky130_fd_sc_hd__nand2_1 _33565_ (.A(_10607_),
    .B(_10624_),
    .Y(_11217_));
 sky130_fd_sc_hd__nand2_4 _33566_ (.A(_11217_),
    .B(_10621_),
    .Y(_11218_));
 sky130_fd_sc_hd__nand3_2 _33567_ (.A(_11210_),
    .B(_11197_),
    .C(_11195_),
    .Y(_11219_));
 sky130_fd_sc_hd__nand3_4 _33568_ (.A(_11216_),
    .B(_11218_),
    .C(_11219_),
    .Y(_11220_));
 sky130_fd_sc_hd__a21o_2 _33569_ (.A1(_10605_),
    .A2(_10603_),
    .B1(_10595_),
    .X(_11221_));
 sky130_fd_sc_hd__a21oi_4 _33570_ (.A1(_11215_),
    .A2(_11220_),
    .B1(_11221_),
    .Y(_11222_));
 sky130_fd_sc_hd__and3_2 _33571_ (.A(_11215_),
    .B(_11220_),
    .C(_11221_),
    .X(_11223_));
 sky130_fd_sc_hd__buf_4 _33572_ (.A(_08787_),
    .X(_11224_));
 sky130_fd_sc_hd__a22oi_4 _33573_ (.A1(_05452_),
    .A2(_09365_),
    .B1(_06505_),
    .B2(_11224_),
    .Y(_11225_));
 sky130_fd_sc_hd__nand3_4 _33574_ (.A(_05587_),
    .B(_06835_),
    .C(_09075_),
    .Y(_11226_));
 sky130_fd_sc_hd__nor2_4 _33575_ (.A(_10652_),
    .B(_11226_),
    .Y(_11227_));
 sky130_fd_sc_hd__buf_4 _33576_ (.A(_19847_),
    .X(_11228_));
 sky130_fd_sc_hd__nand2_2 _33577_ (.A(_05699_),
    .B(_11228_),
    .Y(_11229_));
 sky130_fd_sc_hd__o21ai_2 _33578_ (.A1(_11225_),
    .A2(_11227_),
    .B1(_11229_),
    .Y(_11230_));
 sky130_vsdinv _33579_ (.A(_11229_),
    .Y(_11231_));
 sky130_fd_sc_hd__buf_4 _33580_ (.A(\pcpi_mul.rs1[24] ),
    .X(_11232_));
 sky130_fd_sc_hd__a22o_2 _33581_ (.A1(_05452_),
    .A2(_11232_),
    .B1(_05405_),
    .B2(_09823_),
    .X(_11233_));
 sky130_fd_sc_hd__o211ai_2 _33582_ (.A1(_09929_),
    .A2(_11226_),
    .B1(_11231_),
    .C1(_11233_),
    .Y(_11234_));
 sky130_fd_sc_hd__o21ai_2 _33583_ (.A1(_10743_),
    .A2(_10739_),
    .B1(_10746_),
    .Y(_11235_));
 sky130_fd_sc_hd__nand3_4 _33584_ (.A(_11230_),
    .B(_11234_),
    .C(_11235_),
    .Y(_11236_));
 sky130_fd_sc_hd__a31oi_4 _33585_ (.A1(_10747_),
    .A2(net456),
    .A3(_19864_),
    .B1(_10742_),
    .Y(_11237_));
 sky130_fd_sc_hd__o21ai_2 _33586_ (.A1(_11225_),
    .A2(_11227_),
    .B1(_11231_),
    .Y(_11238_));
 sky130_fd_sc_hd__o211ai_2 _33587_ (.A1(_10652_),
    .A2(_11226_),
    .B1(_11229_),
    .C1(_11233_),
    .Y(_11239_));
 sky130_fd_sc_hd__nand3_4 _33588_ (.A(_11237_),
    .B(_11238_),
    .C(_11239_),
    .Y(_11240_));
 sky130_fd_sc_hd__nor2_8 _33589_ (.A(_10648_),
    .B(_10641_),
    .Y(_11241_));
 sky130_fd_sc_hd__o2bb2ai_4 _33590_ (.A1_N(_11236_),
    .A2_N(_11240_),
    .B1(_10647_),
    .B2(_11241_),
    .Y(_11242_));
 sky130_fd_sc_hd__nor2_4 _33591_ (.A(_10647_),
    .B(_11241_),
    .Y(_11243_));
 sky130_fd_sc_hd__nand3_4 _33592_ (.A(_11240_),
    .B(_11236_),
    .C(_11243_),
    .Y(_11244_));
 sky130_fd_sc_hd__nand2_4 _33593_ (.A(_10750_),
    .B(_10751_),
    .Y(_11245_));
 sky130_fd_sc_hd__a21oi_4 _33594_ (.A1(_11242_),
    .A2(_11244_),
    .B1(_11245_),
    .Y(_11246_));
 sky130_vsdinv _33595_ (.A(_11236_),
    .Y(_11247_));
 sky130_fd_sc_hd__nand2_1 _33596_ (.A(_11240_),
    .B(_11243_),
    .Y(_11248_));
 sky130_fd_sc_hd__o211a_1 _33597_ (.A1(_11247_),
    .A2(_11248_),
    .B1(_11242_),
    .C1(_11245_),
    .X(_11249_));
 sky130_fd_sc_hd__nand2_1 _33598_ (.A(_10656_),
    .B(_10658_),
    .Y(_11250_));
 sky130_fd_sc_hd__nand2_4 _33599_ (.A(_11250_),
    .B(_10650_),
    .Y(_11251_));
 sky130_fd_sc_hd__o21ai_4 _33600_ (.A1(_11246_),
    .A2(_11249_),
    .B1(_11251_),
    .Y(_11252_));
 sky130_fd_sc_hd__a21o_1 _33601_ (.A1(_11242_),
    .A2(_11244_),
    .B1(_11245_),
    .X(_11253_));
 sky130_fd_sc_hd__nand3_4 _33602_ (.A(_11245_),
    .B(_11242_),
    .C(_11244_),
    .Y(_11254_));
 sky130_fd_sc_hd__nand3b_4 _33603_ (.A_N(_11251_),
    .B(_11253_),
    .C(_11254_),
    .Y(_11255_));
 sky130_fd_sc_hd__o21ai_4 _33604_ (.A1(_10673_),
    .A2(_10674_),
    .B1(_10670_),
    .Y(_11256_));
 sky130_fd_sc_hd__a21oi_4 _33605_ (.A1(_11252_),
    .A2(_11255_),
    .B1(_11256_),
    .Y(_11257_));
 sky130_fd_sc_hd__o211a_1 _33606_ (.A1(_10675_),
    .A2(_10680_),
    .B1(_11255_),
    .C1(_11252_),
    .X(_11258_));
 sky130_fd_sc_hd__o22ai_4 _33607_ (.A1(_11222_),
    .A2(_11223_),
    .B1(_11257_),
    .B2(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__a21o_1 _33608_ (.A1(_11252_),
    .A2(_11255_),
    .B1(_11256_),
    .X(_11260_));
 sky130_fd_sc_hd__nor2_2 _33609_ (.A(_11222_),
    .B(_11223_),
    .Y(_11261_));
 sky130_fd_sc_hd__nand3_4 _33610_ (.A(_11252_),
    .B(_11256_),
    .C(_11255_),
    .Y(_11262_));
 sky130_fd_sc_hd__nand3_4 _33611_ (.A(_11260_),
    .B(_11261_),
    .C(_11262_),
    .Y(_11263_));
 sky130_vsdinv _33612_ (.A(_10764_),
    .Y(_11264_));
 sky130_fd_sc_hd__nand2_1 _33613_ (.A(_10757_),
    .B(_10758_),
    .Y(_11265_));
 sky130_fd_sc_hd__o2bb2ai_4 _33614_ (.A1_N(_10771_),
    .A2_N(_10773_),
    .B1(_11264_),
    .B2(_11265_),
    .Y(_11266_));
 sky130_fd_sc_hd__a21oi_2 _33615_ (.A1(_11259_),
    .A2(_11263_),
    .B1(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__nand2_1 _33616_ (.A(_11261_),
    .B(_11262_),
    .Y(_11268_));
 sky130_fd_sc_hd__o211a_1 _33617_ (.A1(_11257_),
    .A2(_11268_),
    .B1(_11266_),
    .C1(_11259_),
    .X(_11269_));
 sky130_fd_sc_hd__a21bo_4 _33618_ (.A1(_10678_),
    .A2(_10685_),
    .B1_N(_10682_),
    .X(_11270_));
 sky130_fd_sc_hd__o21bai_4 _33619_ (.A1(_11267_),
    .A2(_11269_),
    .B1_N(_11270_),
    .Y(_11271_));
 sky130_fd_sc_hd__a21o_1 _33620_ (.A1(_11259_),
    .A2(_11263_),
    .B1(_11266_),
    .X(_11272_));
 sky130_fd_sc_hd__nand3_4 _33621_ (.A(_11259_),
    .B(_11266_),
    .C(_11263_),
    .Y(_11273_));
 sky130_fd_sc_hd__nand3_4 _33622_ (.A(_11272_),
    .B(_11273_),
    .C(_11270_),
    .Y(_11274_));
 sky130_fd_sc_hd__and2_4 _33623_ (.A(_11271_),
    .B(_11274_),
    .X(_11275_));
 sky130_fd_sc_hd__nand2_1 _33624_ (.A(_11177_),
    .B(_11275_),
    .Y(_11276_));
 sky130_fd_sc_hd__a31oi_4 _33625_ (.A1(_10910_),
    .A2(_10916_),
    .A3(_10918_),
    .B1(_10901_),
    .Y(_11277_));
 sky130_fd_sc_hd__nand2_8 _33626_ (.A(_11271_),
    .B(_11274_),
    .Y(_11278_));
 sky130_fd_sc_hd__nand3_2 _33627_ (.A(_11278_),
    .B(_11170_),
    .C(_11176_),
    .Y(_11279_));
 sky130_fd_sc_hd__nand3_4 _33628_ (.A(_11276_),
    .B(_11277_),
    .C(_11279_),
    .Y(_11280_));
 sky130_fd_sc_hd__nand2_1 _33629_ (.A(_11177_),
    .B(_11278_),
    .Y(_11281_));
 sky130_fd_sc_hd__nand3_4 _33630_ (.A(_11275_),
    .B(_11170_),
    .C(_11176_),
    .Y(_11282_));
 sky130_fd_sc_hd__nand3_4 _33631_ (.A(_10910_),
    .B(_10916_),
    .C(_10918_),
    .Y(_11283_));
 sky130_fd_sc_hd__nand2_1 _33632_ (.A(_11283_),
    .B(_10903_),
    .Y(_11284_));
 sky130_fd_sc_hd__nand3_4 _33633_ (.A(_11281_),
    .B(_11282_),
    .C(_11284_),
    .Y(_11285_));
 sky130_fd_sc_hd__nand2_2 _33634_ (.A(_10639_),
    .B(_10629_),
    .Y(_11286_));
 sky130_fd_sc_hd__a21o_2 _33635_ (.A1(_10698_),
    .A2(_10688_),
    .B1(_11286_),
    .X(_11287_));
 sky130_fd_sc_hd__nand3_4 _33636_ (.A(_10698_),
    .B(_10688_),
    .C(_11286_),
    .Y(_11288_));
 sky130_fd_sc_hd__nand3_4 _33637_ (.A(_11287_),
    .B(_18476_),
    .C(_11288_),
    .Y(_11289_));
 sky130_vsdinv _33638_ (.A(_11289_),
    .Y(_11290_));
 sky130_fd_sc_hd__nand2_1 _33639_ (.A(_11287_),
    .B(_11288_),
    .Y(_11291_));
 sky130_fd_sc_hd__buf_4 _33640_ (.A(_11080_),
    .X(_11292_));
 sky130_fd_sc_hd__clkbuf_4 _33641_ (.A(_11292_),
    .X(_11293_));
 sky130_fd_sc_hd__clkbuf_4 _33642_ (.A(_11293_),
    .X(_11294_));
 sky130_fd_sc_hd__nand2_2 _33643_ (.A(_11291_),
    .B(_11294_),
    .Y(_11295_));
 sky130_vsdinv _33644_ (.A(_11295_),
    .Y(_11296_));
 sky130_fd_sc_hd__o2bb2ai_2 _33645_ (.A1_N(_11280_),
    .A2_N(_11285_),
    .B1(_11290_),
    .B2(_11296_),
    .Y(_11297_));
 sky130_fd_sc_hd__nand2_4 _33646_ (.A(_11295_),
    .B(_11289_),
    .Y(_11298_));
 sky130_fd_sc_hd__nand3b_2 _33647_ (.A_N(_11298_),
    .B(_11280_),
    .C(_11285_),
    .Y(_11299_));
 sky130_fd_sc_hd__a21boi_2 _33648_ (.A1(_10936_),
    .A2(_10914_),
    .B1_N(_10924_),
    .Y(_11300_));
 sky130_fd_sc_hd__nand3_4 _33649_ (.A(_11297_),
    .B(_11299_),
    .C(_11300_),
    .Y(_11301_));
 sky130_fd_sc_hd__a21o_1 _33650_ (.A1(_11285_),
    .A2(_11280_),
    .B1(_11298_),
    .X(_11302_));
 sky130_fd_sc_hd__a21bo_1 _33651_ (.A1(_10914_),
    .A2(_10936_),
    .B1_N(_10924_),
    .X(_11303_));
 sky130_fd_sc_hd__nand3_2 _33652_ (.A(_11285_),
    .B(_11280_),
    .C(_11298_),
    .Y(_11304_));
 sky130_fd_sc_hd__nand3_4 _33653_ (.A(_11302_),
    .B(_11303_),
    .C(_11304_),
    .Y(_11305_));
 sky130_fd_sc_hd__o2bb2ai_2 _33654_ (.A1_N(_11301_),
    .A2_N(_11305_),
    .B1(_10926_),
    .B2(_10928_),
    .Y(_11306_));
 sky130_fd_sc_hd__nand3_4 _33655_ (.A(_11305_),
    .B(_11301_),
    .C(_10935_),
    .Y(_11307_));
 sky130_fd_sc_hd__a21bo_1 _33656_ (.A1(_10568_),
    .A2(_10938_),
    .B1_N(_10944_),
    .X(_11308_));
 sky130_fd_sc_hd__a21o_2 _33657_ (.A1(_11306_),
    .A2(_11307_),
    .B1(_11308_),
    .X(_11309_));
 sky130_fd_sc_hd__nand3_4 _33658_ (.A(_11306_),
    .B(_11308_),
    .C(_11307_),
    .Y(_11310_));
 sky130_fd_sc_hd__nand2_4 _33659_ (.A(_11309_),
    .B(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__o2111a_1 _33660_ (.A1(_10586_),
    .A2(_10587_),
    .B1(_09917_),
    .C1(_10240_),
    .D1(_10237_),
    .X(_11312_));
 sky130_fd_sc_hd__nand3_4 _33661_ (.A(_11312_),
    .B(_10585_),
    .C(_10953_),
    .Y(_11313_));
 sky130_fd_sc_hd__nor2_8 _33662_ (.A(_09919_),
    .B(_11313_),
    .Y(_11314_));
 sky130_fd_sc_hd__o2111ai_4 _33663_ (.A1(_06578_),
    .A2(_06393_),
    .B1(_08438_),
    .C1(_06583_),
    .D1(_11314_),
    .Y(_11315_));
 sky130_fd_sc_hd__nand2_1 _33664_ (.A(_08723_),
    .B(_11314_),
    .Y(_11316_));
 sky130_vsdinv _33665_ (.A(_10945_),
    .Y(_11317_));
 sky130_fd_sc_hd__nand2_2 _33666_ (.A(_10951_),
    .B(_10950_),
    .Y(_11318_));
 sky130_fd_sc_hd__nand3_4 _33667_ (.A(_10581_),
    .B(_10578_),
    .C(_10579_),
    .Y(_11319_));
 sky130_fd_sc_hd__a21o_1 _33668_ (.A1(_10578_),
    .A2(_10579_),
    .B1(_10581_),
    .X(_11320_));
 sky130_fd_sc_hd__a21o_1 _33669_ (.A1(_10950_),
    .A2(_10945_),
    .B1(_10951_),
    .X(_11321_));
 sky130_fd_sc_hd__o2111ai_4 _33670_ (.A1(_11317_),
    .A2(_11318_),
    .B1(_11319_),
    .C1(_11320_),
    .D1(_11321_),
    .Y(_11322_));
 sky130_fd_sc_hd__nor2_2 _33671_ (.A(_10588_),
    .B(_11322_),
    .Y(_11323_));
 sky130_fd_sc_hd__o22a_1 _33672_ (.A1(_11317_),
    .A2(_11318_),
    .B1(_11319_),
    .B2(_10952_),
    .X(_11324_));
 sky130_fd_sc_hd__o21ai_2 _33673_ (.A1(_10589_),
    .A2(_11322_),
    .B1(_11324_),
    .Y(_11325_));
 sky130_fd_sc_hd__a21oi_4 _33674_ (.A1(_09924_),
    .A2(_11323_),
    .B1(_11325_),
    .Y(_11326_));
 sky130_fd_sc_hd__nand3_4 _33675_ (.A(_11315_),
    .B(_11316_),
    .C(_11326_),
    .Y(_11327_));
 sky130_fd_sc_hd__xnor2_2 _33676_ (.A(_11311_),
    .B(net409),
    .Y(_02651_));
 sky130_fd_sc_hd__o21ai_4 _33677_ (.A1(_11174_),
    .A2(_11158_),
    .B1(_11165_),
    .Y(_11328_));
 sky130_fd_sc_hd__nor2_1 _33678_ (.A(_11082_),
    .B(_11077_),
    .Y(_11329_));
 sky130_fd_sc_hd__a21oi_2 _33679_ (.A1(_11329_),
    .A2(_11087_),
    .B1(_11085_),
    .Y(_11330_));
 sky130_fd_sc_hd__a21o_1 _33680_ (.A1(_11089_),
    .A2(_11105_),
    .B1(_11330_),
    .X(_11331_));
 sky130_fd_sc_hd__nand3_4 _33681_ (.A(_11075_),
    .B(_11078_),
    .C(_19926_),
    .Y(_11332_));
 sky130_fd_sc_hd__nor2_4 _33682_ (.A(_05281_),
    .B(_11332_),
    .Y(_11333_));
 sky130_fd_sc_hd__a22oi_4 _33683_ (.A1(_10830_),
    .A2(_05127_),
    .B1(_05106_),
    .B2(_11080_),
    .Y(_11334_));
 sky130_fd_sc_hd__nand2_4 _33684_ (.A(_10827_),
    .B(_05263_),
    .Y(_11335_));
 sky130_fd_sc_hd__o21ai_2 _33685_ (.A1(_11333_),
    .A2(_11334_),
    .B1(_11335_),
    .Y(_11336_));
 sky130_vsdinv _33686_ (.A(_11335_),
    .Y(_11337_));
 sky130_vsdinv _33687_ (.A(_11078_),
    .Y(_11338_));
 sky130_fd_sc_hd__o22ai_4 _33688_ (.A1(_05281_),
    .A2(_18473_),
    .B1(_11338_),
    .B2(_05150_),
    .Y(_11339_));
 sky130_fd_sc_hd__o211ai_4 _33689_ (.A1(_05123_),
    .A2(_11332_),
    .B1(_11337_),
    .C1(_11339_),
    .Y(_11340_));
 sky130_fd_sc_hd__o22ai_4 _33690_ (.A1(_05213_),
    .A2(_11076_),
    .B1(_11082_),
    .B2(_11081_),
    .Y(_11341_));
 sky130_fd_sc_hd__nand3_4 _33691_ (.A(_11336_),
    .B(_11340_),
    .C(_11341_),
    .Y(_11342_));
 sky130_fd_sc_hd__o21ai_2 _33692_ (.A1(_11333_),
    .A2(_11334_),
    .B1(_11337_),
    .Y(_11343_));
 sky130_fd_sc_hd__nand3b_4 _33693_ (.A_N(_11333_),
    .B(_11339_),
    .C(_11335_),
    .Y(_11344_));
 sky130_fd_sc_hd__a21oi_2 _33694_ (.A1(_11087_),
    .A2(_11083_),
    .B1(_11077_),
    .Y(_11345_));
 sky130_fd_sc_hd__nand3_4 _33695_ (.A(_11343_),
    .B(_11344_),
    .C(_11345_),
    .Y(_11346_));
 sky130_fd_sc_hd__nand2_4 _33696_ (.A(_19591_),
    .B(_05486_),
    .Y(_11347_));
 sky130_fd_sc_hd__buf_6 _33697_ (.A(_10835_),
    .X(_11348_));
 sky130_fd_sc_hd__a22oi_4 _33698_ (.A1(_11348_),
    .A2(_19920_),
    .B1(net494),
    .B2(_05268_),
    .Y(_11349_));
 sky130_fd_sc_hd__nand2_1 _33699_ (.A(_10835_),
    .B(_19919_),
    .Y(_11350_));
 sky130_fd_sc_hd__nand2_1 _33700_ (.A(_19586_),
    .B(_19916_),
    .Y(_11351_));
 sky130_fd_sc_hd__nor2_1 _33701_ (.A(_11350_),
    .B(_11351_),
    .Y(_11352_));
 sky130_fd_sc_hd__buf_2 _33702_ (.A(_11352_),
    .X(_11353_));
 sky130_fd_sc_hd__nor3_2 _33703_ (.A(_11347_),
    .B(_11349_),
    .C(_11353_),
    .Y(_11354_));
 sky130_vsdinv _33704_ (.A(_11347_),
    .Y(_11355_));
 sky130_fd_sc_hd__nor2_1 _33705_ (.A(_11349_),
    .B(_11353_),
    .Y(_11356_));
 sky130_fd_sc_hd__nor2_1 _33706_ (.A(_11355_),
    .B(_11356_),
    .Y(_11357_));
 sky130_fd_sc_hd__o2bb2ai_1 _33707_ (.A1_N(_11342_),
    .A2_N(_11346_),
    .B1(_11354_),
    .B2(_11357_),
    .Y(_11358_));
 sky130_fd_sc_hd__nand2_1 _33708_ (.A(_11350_),
    .B(_11351_),
    .Y(_11359_));
 sky130_fd_sc_hd__nand3b_2 _33709_ (.A_N(_11352_),
    .B(_11359_),
    .C(_11347_),
    .Y(_11360_));
 sky130_fd_sc_hd__o21ai_2 _33710_ (.A1(_11349_),
    .A2(_11353_),
    .B1(_11355_),
    .Y(_11361_));
 sky130_fd_sc_hd__nand2_2 _33711_ (.A(_11360_),
    .B(_11361_),
    .Y(_11362_));
 sky130_fd_sc_hd__nand3_2 _33712_ (.A(_11346_),
    .B(_11342_),
    .C(_11362_),
    .Y(_11363_));
 sky130_fd_sc_hd__nand3_4 _33713_ (.A(_11331_),
    .B(_11358_),
    .C(_11363_),
    .Y(_11364_));
 sky130_vsdinv _33714_ (.A(_11361_),
    .Y(_11365_));
 sky130_vsdinv _33715_ (.A(_11360_),
    .Y(_11366_));
 sky130_fd_sc_hd__o2bb2ai_1 _33716_ (.A1_N(_11342_),
    .A2_N(_11346_),
    .B1(_11365_),
    .B2(_11366_),
    .Y(_11367_));
 sky130_fd_sc_hd__a21oi_2 _33717_ (.A1(_11089_),
    .A2(_11105_),
    .B1(_11330_),
    .Y(_11368_));
 sky130_fd_sc_hd__nand3b_2 _33718_ (.A_N(_11362_),
    .B(_11342_),
    .C(_11346_),
    .Y(_11369_));
 sky130_fd_sc_hd__nand3_4 _33719_ (.A(_11367_),
    .B(_11368_),
    .C(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__nand2_1 _33720_ (.A(_11364_),
    .B(_11370_),
    .Y(_11371_));
 sky130_fd_sc_hd__o21a_2 _33721_ (.A1(_11114_),
    .A2(_11112_),
    .B1(_11119_),
    .X(_11372_));
 sky130_fd_sc_hd__nand2_2 _33722_ (.A(_10256_),
    .B(_08198_),
    .Y(_11373_));
 sky130_fd_sc_hd__nand2_2 _33723_ (.A(_08946_),
    .B(_05672_),
    .Y(_11374_));
 sky130_fd_sc_hd__nor2_2 _33724_ (.A(_11373_),
    .B(_11374_),
    .Y(_11375_));
 sky130_fd_sc_hd__nor2_4 _33725_ (.A(_08578_),
    .B(_05802_),
    .Y(_11376_));
 sky130_fd_sc_hd__nand2_2 _33726_ (.A(_11373_),
    .B(_11374_),
    .Y(_11377_));
 sky130_fd_sc_hd__nand3b_4 _33727_ (.A_N(_11375_),
    .B(_11376_),
    .C(_11377_),
    .Y(_11378_));
 sky130_fd_sc_hd__buf_6 _33728_ (.A(_08946_),
    .X(_11379_));
 sky130_fd_sc_hd__a21o_1 _33729_ (.A1(_11379_),
    .A2(_05808_),
    .B1(_11373_),
    .X(_11380_));
 sky130_fd_sc_hd__a21o_1 _33730_ (.A1(_19597_),
    .A2(_05671_),
    .B1(_11374_),
    .X(_11381_));
 sky130_fd_sc_hd__o211ai_4 _33731_ (.A1(_08579_),
    .A2(_05981_),
    .B1(_11380_),
    .C1(_11381_),
    .Y(_11382_));
 sky130_fd_sc_hd__a21o_2 _33732_ (.A1(_11100_),
    .A2(_11098_),
    .B1(_11096_),
    .X(_11383_));
 sky130_fd_sc_hd__a21oi_4 _33733_ (.A1(_11378_),
    .A2(_11382_),
    .B1(_11383_),
    .Y(_11384_));
 sky130_fd_sc_hd__nor2_2 _33734_ (.A(_11372_),
    .B(_11384_),
    .Y(_11385_));
 sky130_fd_sc_hd__nand3_4 _33735_ (.A(_11383_),
    .B(_11378_),
    .C(_11382_),
    .Y(_11386_));
 sky130_fd_sc_hd__nor2_1 _33736_ (.A(_11098_),
    .B(_11096_),
    .Y(_11387_));
 sky130_fd_sc_hd__o2bb2ai_1 _33737_ (.A1_N(_11382_),
    .A2_N(_11378_),
    .B1(_11093_),
    .B2(_11387_),
    .Y(_11388_));
 sky130_fd_sc_hd__o21ai_2 _33738_ (.A1(_11114_),
    .A2(_11112_),
    .B1(_11119_),
    .Y(_11389_));
 sky130_fd_sc_hd__a21oi_2 _33739_ (.A1(_11388_),
    .A2(_11386_),
    .B1(_11389_),
    .Y(_11390_));
 sky130_fd_sc_hd__a21oi_4 _33740_ (.A1(_11385_),
    .A2(_11386_),
    .B1(_11390_),
    .Y(_11391_));
 sky130_fd_sc_hd__nand2_1 _33741_ (.A(_11371_),
    .B(_11391_),
    .Y(_11392_));
 sky130_fd_sc_hd__a21boi_4 _33742_ (.A1(_11131_),
    .A2(_11110_),
    .B1_N(_11107_),
    .Y(_11393_));
 sky130_fd_sc_hd__nand2_1 _33743_ (.A(_11385_),
    .B(_11386_),
    .Y(_11394_));
 sky130_fd_sc_hd__a21o_1 _33744_ (.A1(_11388_),
    .A2(_11386_),
    .B1(_11389_),
    .X(_11395_));
 sky130_fd_sc_hd__nand2_1 _33745_ (.A(_11394_),
    .B(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__nand3_2 _33746_ (.A(_11396_),
    .B(_11370_),
    .C(_11364_),
    .Y(_11397_));
 sky130_fd_sc_hd__nand3_4 _33747_ (.A(_11392_),
    .B(_11393_),
    .C(_11397_),
    .Y(_11398_));
 sky130_fd_sc_hd__nand2_2 _33748_ (.A(_11371_),
    .B(_11396_),
    .Y(_11399_));
 sky130_fd_sc_hd__o2bb2ai_2 _33749_ (.A1_N(_11131_),
    .A2_N(_11110_),
    .B1(_11140_),
    .B2(_11144_),
    .Y(_11400_));
 sky130_fd_sc_hd__nand3_4 _33750_ (.A(_11391_),
    .B(_11370_),
    .C(_11364_),
    .Y(_11401_));
 sky130_fd_sc_hd__nand3_4 _33751_ (.A(_11399_),
    .B(_11400_),
    .C(_11401_),
    .Y(_11402_));
 sky130_fd_sc_hd__nand2_1 _33752_ (.A(_11398_),
    .B(_11402_),
    .Y(_11403_));
 sky130_fd_sc_hd__a22oi_4 _33753_ (.A1(_10073_),
    .A2(_07789_),
    .B1(_10066_),
    .B2(_19898_),
    .Y(_11404_));
 sky130_fd_sc_hd__nand3_4 _33754_ (.A(_08539_),
    .B(_08154_),
    .C(_06259_),
    .Y(_11405_));
 sky130_fd_sc_hd__nor2_4 _33755_ (.A(_05787_),
    .B(_11405_),
    .Y(_11406_));
 sky130_fd_sc_hd__nand2_4 _33756_ (.A(_19615_),
    .B(_19893_),
    .Y(_11407_));
 sky130_fd_sc_hd__o21ai_2 _33757_ (.A1(_11404_),
    .A2(_11406_),
    .B1(_11407_),
    .Y(_11408_));
 sky130_fd_sc_hd__o22ai_4 _33758_ (.A1(net442),
    .A2(_10791_),
    .B1(_11040_),
    .B2(_11044_),
    .Y(_11409_));
 sky130_vsdinv _33759_ (.A(_11407_),
    .Y(_11410_));
 sky130_fd_sc_hd__a22o_1 _33760_ (.A1(_10073_),
    .A2(_07789_),
    .B1(_09680_),
    .B2(_06657_),
    .X(_11411_));
 sky130_fd_sc_hd__o211ai_2 _33761_ (.A1(_07102_),
    .A2(_11405_),
    .B1(_11410_),
    .C1(_11411_),
    .Y(_11412_));
 sky130_fd_sc_hd__nand3_4 _33762_ (.A(_11408_),
    .B(_11409_),
    .C(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__o21ai_2 _33763_ (.A1(_11404_),
    .A2(_11406_),
    .B1(_11410_),
    .Y(_11414_));
 sky130_fd_sc_hd__a21oi_2 _33764_ (.A1(_11042_),
    .A2(_11041_),
    .B1(_11045_),
    .Y(_11415_));
 sky130_fd_sc_hd__o211ai_2 _33765_ (.A1(_07102_),
    .A2(_11405_),
    .B1(_11407_),
    .C1(_11411_),
    .Y(_11416_));
 sky130_fd_sc_hd__nand3_4 _33766_ (.A(_11414_),
    .B(_11415_),
    .C(_11416_),
    .Y(_11417_));
 sky130_fd_sc_hd__a22oi_4 _33767_ (.A1(_07978_),
    .A2(_07072_),
    .B1(_19625_),
    .B2(_07330_),
    .Y(_11418_));
 sky130_fd_sc_hd__nand2_2 _33768_ (.A(_07822_),
    .B(_06779_),
    .Y(_11419_));
 sky130_fd_sc_hd__nand2_2 _33769_ (.A(_07827_),
    .B(_06267_),
    .Y(_11420_));
 sky130_fd_sc_hd__nor2_2 _33770_ (.A(_11419_),
    .B(_11420_),
    .Y(_11421_));
 sky130_fd_sc_hd__nand2_2 _33771_ (.A(_10364_),
    .B(_06641_),
    .Y(_11422_));
 sky130_fd_sc_hd__o21a_1 _33772_ (.A1(_11418_),
    .A2(_11421_),
    .B1(_11422_),
    .X(_11423_));
 sky130_fd_sc_hd__nor3_4 _33773_ (.A(_11422_),
    .B(_11418_),
    .C(_11421_),
    .Y(_11424_));
 sky130_fd_sc_hd__o2bb2ai_2 _33774_ (.A1_N(_11413_),
    .A2_N(_11417_),
    .B1(_11423_),
    .B2(_11424_),
    .Y(_11425_));
 sky130_fd_sc_hd__o21ai_2 _33775_ (.A1(_11125_),
    .A2(_11127_),
    .B1(_11123_),
    .Y(_11426_));
 sky130_fd_sc_hd__nor2_2 _33776_ (.A(_11424_),
    .B(_11423_),
    .Y(_11427_));
 sky130_fd_sc_hd__nand3_4 _33777_ (.A(_11427_),
    .B(_11417_),
    .C(_11413_),
    .Y(_11428_));
 sky130_fd_sc_hd__and3_4 _33778_ (.A(_11425_),
    .B(_11426_),
    .C(_11428_),
    .X(_11429_));
 sky130_fd_sc_hd__a21o_1 _33779_ (.A1(_11425_),
    .A2(_11428_),
    .B1(_11426_),
    .X(_11430_));
 sky130_fd_sc_hd__nand2_2 _33780_ (.A(_11148_),
    .B(_11047_),
    .Y(_11431_));
 sky130_fd_sc_hd__nand2_2 _33781_ (.A(_11430_),
    .B(_11431_),
    .Y(_11432_));
 sky130_fd_sc_hd__a21oi_1 _33782_ (.A1(_11425_),
    .A2(_11428_),
    .B1(_11426_),
    .Y(_11433_));
 sky130_fd_sc_hd__o21bai_2 _33783_ (.A1(_11433_),
    .A2(_11429_),
    .B1_N(_11431_),
    .Y(_11434_));
 sky130_fd_sc_hd__o21ai_4 _33784_ (.A1(_11429_),
    .A2(_11432_),
    .B1(_11434_),
    .Y(_11435_));
 sky130_fd_sc_hd__nand2_2 _33785_ (.A(_11403_),
    .B(_11435_),
    .Y(_11436_));
 sky130_vsdinv _33786_ (.A(_10789_),
    .Y(_11437_));
 sky130_fd_sc_hd__and3_1 _33787_ (.A(_10804_),
    .B(_10801_),
    .C(_10799_),
    .X(_11438_));
 sky130_fd_sc_hd__o22ai_2 _33788_ (.A1(_11437_),
    .A2(_11438_),
    .B1(_11147_),
    .B2(_11150_),
    .Y(_11439_));
 sky130_fd_sc_hd__nand2_2 _33789_ (.A(_11439_),
    .B(_11073_),
    .Y(_11440_));
 sky130_fd_sc_hd__o22ai_4 _33790_ (.A1(_11145_),
    .A2(_11162_),
    .B1(_11440_),
    .B2(_11135_),
    .Y(_11441_));
 sky130_fd_sc_hd__o21a_1 _33791_ (.A1(_11429_),
    .A2(_11432_),
    .B1(_11434_),
    .X(_11442_));
 sky130_fd_sc_hd__nand3_4 _33792_ (.A(_11442_),
    .B(_11398_),
    .C(_11402_),
    .Y(_11443_));
 sky130_fd_sc_hd__nand3_4 _33793_ (.A(_11436_),
    .B(_11441_),
    .C(_11443_),
    .Y(_11444_));
 sky130_fd_sc_hd__a21oi_4 _33794_ (.A1(_11146_),
    .A2(_11154_),
    .B1(_11137_),
    .Y(_11445_));
 sky130_fd_sc_hd__nand2_1 _33795_ (.A(_11403_),
    .B(_11442_),
    .Y(_11446_));
 sky130_fd_sc_hd__nand3_2 _33796_ (.A(_11435_),
    .B(_11398_),
    .C(_11402_),
    .Y(_11447_));
 sky130_fd_sc_hd__nand3_4 _33797_ (.A(_11445_),
    .B(_11446_),
    .C(_11447_),
    .Y(_11448_));
 sky130_fd_sc_hd__a21oi_4 _33798_ (.A1(_11019_),
    .A2(_11032_),
    .B1(_11017_),
    .Y(_11449_));
 sky130_fd_sc_hd__nand3_4 _33799_ (.A(_19632_),
    .B(_08616_),
    .C(_19881_),
    .Y(_11450_));
 sky130_fd_sc_hd__nor2_4 _33800_ (.A(_08447_),
    .B(_11450_),
    .Y(_11451_));
 sky130_fd_sc_hd__a22o_2 _33801_ (.A1(_10990_),
    .A2(_06804_),
    .B1(_19637_),
    .B2(_07344_),
    .X(_11452_));
 sky130_fd_sc_hd__nand2_2 _33802_ (.A(_07435_),
    .B(_19874_),
    .Y(_11453_));
 sky130_fd_sc_hd__nand3b_4 _33803_ (.A_N(_11451_),
    .B(_11452_),
    .C(_11453_),
    .Y(_11454_));
 sky130_fd_sc_hd__nand2_1 _33804_ (.A(_11056_),
    .B(_11057_),
    .Y(_11455_));
 sky130_fd_sc_hd__a21oi_2 _33805_ (.A1(_11054_),
    .A2(_11455_),
    .B1(_11058_),
    .Y(_11456_));
 sky130_fd_sc_hd__a22oi_4 _33806_ (.A1(_19633_),
    .A2(_19882_),
    .B1(_19637_),
    .B2(_19879_),
    .Y(_11457_));
 sky130_vsdinv _33807_ (.A(_11453_),
    .Y(_11458_));
 sky130_fd_sc_hd__o21ai_2 _33808_ (.A1(_11457_),
    .A2(_11451_),
    .B1(_11458_),
    .Y(_11459_));
 sky130_fd_sc_hd__nand3_4 _33809_ (.A(_11454_),
    .B(_11456_),
    .C(_11459_),
    .Y(_11460_));
 sky130_fd_sc_hd__nor2_2 _33810_ (.A(_11053_),
    .B(_11055_),
    .Y(_11461_));
 sky130_fd_sc_hd__o211ai_4 _33811_ (.A1(net438),
    .A2(_11450_),
    .B1(_11458_),
    .C1(_11452_),
    .Y(_11462_));
 sky130_fd_sc_hd__o21ai_2 _33812_ (.A1(_11457_),
    .A2(_11451_),
    .B1(_11453_),
    .Y(_11463_));
 sky130_fd_sc_hd__o211ai_4 _33813_ (.A1(_11058_),
    .A2(_11461_),
    .B1(_11462_),
    .C1(_11463_),
    .Y(_11464_));
 sky130_fd_sc_hd__a21o_2 _33814_ (.A1(_11000_),
    .A2(_10996_),
    .B1(_10994_),
    .X(_11465_));
 sky130_fd_sc_hd__a21o_2 _33815_ (.A1(_11460_),
    .A2(_11464_),
    .B1(_11465_),
    .X(_11466_));
 sky130_fd_sc_hd__nand3_4 _33816_ (.A(_11460_),
    .B(_11464_),
    .C(_11465_),
    .Y(_11467_));
 sky130_fd_sc_hd__nand2_4 _33817_ (.A(_11012_),
    .B(_11007_),
    .Y(_11468_));
 sky130_fd_sc_hd__a21oi_4 _33818_ (.A1(_11466_),
    .A2(_11467_),
    .B1(_11468_),
    .Y(_11469_));
 sky130_vsdinv _33819_ (.A(_11007_),
    .Y(_11470_));
 sky130_fd_sc_hd__o21a_1 _33820_ (.A1(_10706_),
    .A2(_11011_),
    .B1(_11002_),
    .X(_11471_));
 sky130_fd_sc_hd__o211a_1 _33821_ (.A1(_11470_),
    .A2(_11471_),
    .B1(_11467_),
    .C1(_11466_),
    .X(_11472_));
 sky130_fd_sc_hd__nand3_4 _33822_ (.A(_06411_),
    .B(_06169_),
    .C(_08062_),
    .Y(_11473_));
 sky130_fd_sc_hd__a22o_2 _33823_ (.A1(_06606_),
    .A2(_19871_),
    .B1(_09439_),
    .B2(_07705_),
    .X(_11474_));
 sky130_fd_sc_hd__o21ai_1 _33824_ (.A1(_10654_),
    .A2(_11473_),
    .B1(_11474_),
    .Y(_11475_));
 sky130_fd_sc_hd__nand2_2 _33825_ (.A(_06349_),
    .B(_08336_),
    .Y(_11476_));
 sky130_fd_sc_hd__nand2_1 _33826_ (.A(_11475_),
    .B(_11476_),
    .Y(_11477_));
 sky130_fd_sc_hd__a21o_1 _33827_ (.A1(_10965_),
    .A2(_10966_),
    .B1(_10962_),
    .X(_11478_));
 sky130_fd_sc_hd__nor2_1 _33828_ (.A(_10654_),
    .B(_11473_),
    .Y(_11479_));
 sky130_vsdinv _33829_ (.A(_11476_),
    .Y(_11480_));
 sky130_fd_sc_hd__nand3b_2 _33830_ (.A_N(_11479_),
    .B(_11474_),
    .C(_11480_),
    .Y(_11481_));
 sky130_fd_sc_hd__nand3_4 _33831_ (.A(_11477_),
    .B(_11478_),
    .C(_11481_),
    .Y(_11482_));
 sky130_vsdinv _33832_ (.A(_11482_),
    .Y(_11483_));
 sky130_fd_sc_hd__a22oi_4 _33833_ (.A1(_06327_),
    .A2(_08332_),
    .B1(_05737_),
    .B2(_09082_),
    .Y(_11484_));
 sky130_fd_sc_hd__and4_2 _33834_ (.A(_06398_),
    .B(_19655_),
    .C(_10459_),
    .D(_10458_),
    .X(_11485_));
 sky130_fd_sc_hd__nor2_1 _33835_ (.A(_11484_),
    .B(_11485_),
    .Y(_11486_));
 sky130_fd_sc_hd__nand2_2 _33836_ (.A(_05732_),
    .B(_09365_),
    .Y(_11487_));
 sky130_fd_sc_hd__nand2_1 _33837_ (.A(_11486_),
    .B(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__o21bai_2 _33838_ (.A1(_11484_),
    .A2(_11485_),
    .B1_N(_11487_),
    .Y(_11489_));
 sky130_fd_sc_hd__nand2_4 _33839_ (.A(_11488_),
    .B(_11489_),
    .Y(_11490_));
 sky130_fd_sc_hd__nand2_1 _33840_ (.A(_11475_),
    .B(_11480_),
    .Y(_11491_));
 sky130_fd_sc_hd__a21oi_2 _33841_ (.A1(_10965_),
    .A2(_10966_),
    .B1(_10962_),
    .Y(_11492_));
 sky130_fd_sc_hd__o211ai_4 _33842_ (.A1(_08080_),
    .A2(_11473_),
    .B1(_11476_),
    .C1(_11474_),
    .Y(_11493_));
 sky130_fd_sc_hd__nand3_4 _33843_ (.A(_11491_),
    .B(_11492_),
    .C(_11493_),
    .Y(_11494_));
 sky130_fd_sc_hd__nand2_4 _33844_ (.A(_11490_),
    .B(_11494_),
    .Y(_11495_));
 sky130_vsdinv _33845_ (.A(_11490_),
    .Y(_11496_));
 sky130_fd_sc_hd__nand2_1 _33846_ (.A(_11482_),
    .B(_11494_),
    .Y(_11497_));
 sky130_fd_sc_hd__nand2_2 _33847_ (.A(_11496_),
    .B(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__o21ai_4 _33848_ (.A1(_11483_),
    .A2(_11495_),
    .B1(_11498_),
    .Y(_11499_));
 sky130_fd_sc_hd__o21ai_2 _33849_ (.A1(_11469_),
    .A2(_11472_),
    .B1(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__a21o_1 _33850_ (.A1(_11466_),
    .A2(_11467_),
    .B1(_11468_),
    .X(_11501_));
 sky130_fd_sc_hd__o21a_1 _33851_ (.A1(_11483_),
    .A2(_11495_),
    .B1(_11498_),
    .X(_11502_));
 sky130_fd_sc_hd__nand3_4 _33852_ (.A(_11468_),
    .B(_11466_),
    .C(_11467_),
    .Y(_11503_));
 sky130_fd_sc_hd__nand3_2 _33853_ (.A(_11501_),
    .B(_11502_),
    .C(_11503_),
    .Y(_11504_));
 sky130_fd_sc_hd__o21ai_2 _33854_ (.A1(_11152_),
    .A2(_11147_),
    .B1(_11069_),
    .Y(_11505_));
 sky130_fd_sc_hd__nand3_4 _33855_ (.A(_11500_),
    .B(_11504_),
    .C(_11505_),
    .Y(_11506_));
 sky130_fd_sc_hd__nor2_2 _33856_ (.A(_11490_),
    .B(_11497_),
    .Y(_11507_));
 sky130_fd_sc_hd__and2_1 _33857_ (.A(_11482_),
    .B(_11494_),
    .X(_11508_));
 sky130_fd_sc_hd__nor2_2 _33858_ (.A(_11496_),
    .B(_11508_),
    .Y(_11509_));
 sky130_fd_sc_hd__o22ai_4 _33859_ (.A1(_11507_),
    .A2(_11509_),
    .B1(_11469_),
    .B2(_11472_),
    .Y(_11510_));
 sky130_fd_sc_hd__nand2_1 _33860_ (.A(_11069_),
    .B(_11152_),
    .Y(_11511_));
 sky130_fd_sc_hd__nand2_4 _33861_ (.A(_11511_),
    .B(_11068_),
    .Y(_11512_));
 sky130_fd_sc_hd__nand3_4 _33862_ (.A(_11501_),
    .B(_11499_),
    .C(_11503_),
    .Y(_11513_));
 sky130_fd_sc_hd__nand3_4 _33863_ (.A(_11510_),
    .B(_11512_),
    .C(_11513_),
    .Y(_11514_));
 sky130_fd_sc_hd__nand2_1 _33864_ (.A(_11506_),
    .B(_11514_),
    .Y(_11515_));
 sky130_fd_sc_hd__nor2_1 _33865_ (.A(_11449_),
    .B(_11515_),
    .Y(_11516_));
 sky130_fd_sc_hd__o21ai_2 _33866_ (.A1(_11024_),
    .A2(_11015_),
    .B1(_11020_),
    .Y(_11517_));
 sky130_fd_sc_hd__a21oi_4 _33867_ (.A1(_11506_),
    .A2(_11514_),
    .B1(_11517_),
    .Y(_11518_));
 sky130_fd_sc_hd__o2bb2ai_2 _33868_ (.A1_N(_11444_),
    .A2_N(_11448_),
    .B1(_11516_),
    .B2(_11518_),
    .Y(_11519_));
 sky130_fd_sc_hd__a31oi_4 _33869_ (.A1(_11510_),
    .A2(_11513_),
    .A3(_11512_),
    .B1(_11449_),
    .Y(_11520_));
 sky130_fd_sc_hd__a21oi_4 _33870_ (.A1(_11506_),
    .A2(_11520_),
    .B1(_11518_),
    .Y(_11521_));
 sky130_fd_sc_hd__nand3_4 _33871_ (.A(_11521_),
    .B(_11448_),
    .C(_11444_),
    .Y(_11522_));
 sky130_fd_sc_hd__nand3_4 _33872_ (.A(_11328_),
    .B(_11519_),
    .C(_11522_),
    .Y(_11523_));
 sky130_fd_sc_hd__nand2_1 _33873_ (.A(_11146_),
    .B(_11155_),
    .Y(_11524_));
 sky130_fd_sc_hd__a22oi_4 _33874_ (.A1(_10880_),
    .A2(_10878_),
    .B1(_11524_),
    .B2(_11440_),
    .Y(_11525_));
 sky130_fd_sc_hd__a22oi_4 _33875_ (.A1(_11156_),
    .A2(_11525_),
    .B1(_11164_),
    .B2(_11168_),
    .Y(_11526_));
 sky130_fd_sc_hd__nand2_1 _33876_ (.A(_11515_),
    .B(_11449_),
    .Y(_11527_));
 sky130_fd_sc_hd__nand2_1 _33877_ (.A(_11520_),
    .B(_11506_),
    .Y(_11528_));
 sky130_fd_sc_hd__nand2_2 _33878_ (.A(_11527_),
    .B(_11528_),
    .Y(_11529_));
 sky130_fd_sc_hd__nand3_2 _33879_ (.A(_11529_),
    .B(_11448_),
    .C(_11444_),
    .Y(_11530_));
 sky130_fd_sc_hd__a21o_1 _33880_ (.A1(_11448_),
    .A2(_11444_),
    .B1(_11529_),
    .X(_11531_));
 sky130_fd_sc_hd__nand3_4 _33881_ (.A(_11526_),
    .B(_11530_),
    .C(_11531_),
    .Y(_11532_));
 sky130_fd_sc_hd__o21a_1 _33882_ (.A1(_11251_),
    .A2(_11246_),
    .B1(_11254_),
    .X(_11533_));
 sky130_vsdinv _33883_ (.A(_11248_),
    .Y(_11534_));
 sky130_fd_sc_hd__a22oi_4 _33884_ (.A1(_05841_),
    .A2(_09362_),
    .B1(_05843_),
    .B2(_09820_),
    .Y(_11535_));
 sky130_vsdinv _33885_ (.A(\pcpi_mul.rs1[25] ),
    .Y(_11536_));
 sky130_fd_sc_hd__clkbuf_8 _33886_ (.A(_11536_),
    .X(_11537_));
 sky130_fd_sc_hd__nand3_4 _33887_ (.A(_06502_),
    .B(_06504_),
    .C(_19848_),
    .Y(_11538_));
 sky130_fd_sc_hd__nor2_8 _33888_ (.A(_11537_),
    .B(_11538_),
    .Y(_11539_));
 sky130_fd_sc_hd__nand2_2 _33889_ (.A(_05699_),
    .B(_09950_),
    .Y(_11540_));
 sky130_vsdinv _33890_ (.A(_11540_),
    .Y(_11541_));
 sky130_fd_sc_hd__o21ai_2 _33891_ (.A1(_11535_),
    .A2(_11539_),
    .B1(_11541_),
    .Y(_11542_));
 sky130_vsdinv _33892_ (.A(_10979_),
    .Y(_11543_));
 sky130_fd_sc_hd__a21oi_2 _33893_ (.A1(_11543_),
    .A2(_10983_),
    .B1(_10978_),
    .Y(_11544_));
 sky130_fd_sc_hd__buf_6 _33894_ (.A(_11536_),
    .X(_11545_));
 sky130_fd_sc_hd__a22o_2 _33895_ (.A1(_05452_),
    .A2(_09362_),
    .B1(_05843_),
    .B2(_09359_),
    .X(_11546_));
 sky130_fd_sc_hd__o211ai_4 _33896_ (.A1(_11545_),
    .A2(_11538_),
    .B1(_11540_),
    .C1(_11546_),
    .Y(_11547_));
 sky130_fd_sc_hd__nand3_4 _33897_ (.A(_11542_),
    .B(_11544_),
    .C(_11547_),
    .Y(_11548_));
 sky130_fd_sc_hd__o21ai_2 _33898_ (.A1(_11535_),
    .A2(_11539_),
    .B1(_11540_),
    .Y(_11549_));
 sky130_fd_sc_hd__o21ai_2 _33899_ (.A1(_10979_),
    .A2(_10975_),
    .B1(_10982_),
    .Y(_11550_));
 sky130_fd_sc_hd__o211ai_4 _33900_ (.A1(_11545_),
    .A2(_11538_),
    .B1(_11541_),
    .C1(_11546_),
    .Y(_11551_));
 sky130_fd_sc_hd__nand3_4 _33901_ (.A(_11549_),
    .B(_11550_),
    .C(_11551_),
    .Y(_11552_));
 sky130_fd_sc_hd__nand2_1 _33902_ (.A(_11548_),
    .B(_11552_),
    .Y(_11553_));
 sky130_fd_sc_hd__a21oi_4 _33903_ (.A1(_11233_),
    .A2(_11231_),
    .B1(_11227_),
    .Y(_11554_));
 sky130_fd_sc_hd__nand2_4 _33904_ (.A(_11553_),
    .B(_11554_),
    .Y(_11555_));
 sky130_fd_sc_hd__nand3b_4 _33905_ (.A_N(_11554_),
    .B(_11548_),
    .C(_11552_),
    .Y(_11556_));
 sky130_fd_sc_hd__nand2_4 _33906_ (.A(_11022_),
    .B(_10968_),
    .Y(_11557_));
 sky130_fd_sc_hd__a21oi_4 _33907_ (.A1(_11555_),
    .A2(_11556_),
    .B1(_11557_),
    .Y(_11558_));
 sky130_fd_sc_hd__a32oi_2 _33908_ (.A1(_10969_),
    .A2(_10970_),
    .A3(_10972_),
    .B1(_10980_),
    .B2(_10984_),
    .Y(_11559_));
 sky130_fd_sc_hd__o211a_2 _33909_ (.A1(_11021_),
    .A2(_11559_),
    .B1(_11556_),
    .C1(_11555_),
    .X(_11560_));
 sky130_fd_sc_hd__o22ai_4 _33910_ (.A1(_11247_),
    .A2(_11534_),
    .B1(_11558_),
    .B2(_11560_),
    .Y(_11561_));
 sky130_fd_sc_hd__a21o_1 _33911_ (.A1(_11555_),
    .A2(_11556_),
    .B1(_11557_),
    .X(_11562_));
 sky130_fd_sc_hd__nand3_4 _33912_ (.A(_11557_),
    .B(_11555_),
    .C(_11556_),
    .Y(_11563_));
 sky130_fd_sc_hd__nor2_4 _33913_ (.A(_11247_),
    .B(_11534_),
    .Y(_11564_));
 sky130_fd_sc_hd__nand3_2 _33914_ (.A(_11562_),
    .B(_11563_),
    .C(_11564_),
    .Y(_11565_));
 sky130_fd_sc_hd__nand3_4 _33915_ (.A(_11533_),
    .B(_11561_),
    .C(_11565_),
    .Y(_11566_));
 sky130_vsdinv _33916_ (.A(_11240_),
    .Y(_11567_));
 sky130_fd_sc_hd__nor2_2 _33917_ (.A(_11243_),
    .B(_11247_),
    .Y(_11568_));
 sky130_fd_sc_hd__o22ai_4 _33918_ (.A1(_11567_),
    .A2(_11568_),
    .B1(_11558_),
    .B2(_11560_),
    .Y(_11569_));
 sky130_fd_sc_hd__nand3b_2 _33919_ (.A_N(_11564_),
    .B(_11562_),
    .C(_11563_),
    .Y(_11570_));
 sky130_fd_sc_hd__o21ai_2 _33920_ (.A1(_11251_),
    .A2(_11246_),
    .B1(_11254_),
    .Y(_11571_));
 sky130_fd_sc_hd__nand3_4 _33921_ (.A(_11569_),
    .B(_11570_),
    .C(_11571_),
    .Y(_11572_));
 sky130_fd_sc_hd__nand2_1 _33922_ (.A(_11566_),
    .B(_11572_),
    .Y(_11573_));
 sky130_fd_sc_hd__buf_6 _33923_ (.A(_10488_),
    .X(_11574_));
 sky130_fd_sc_hd__a22oi_4 _33924_ (.A1(net455),
    .A2(_11574_),
    .B1(_19674_),
    .B2(_19835_),
    .Y(_11575_));
 sky130_fd_sc_hd__nand2_2 _33925_ (.A(_05791_),
    .B(_09946_),
    .Y(_11576_));
 sky130_fd_sc_hd__nand2_2 _33926_ (.A(_05792_),
    .B(_10487_),
    .Y(_11577_));
 sky130_fd_sc_hd__nor2_4 _33927_ (.A(_11576_),
    .B(_11577_),
    .Y(_11578_));
 sky130_fd_sc_hd__buf_2 _33928_ (.A(_11186_),
    .X(_11579_));
 sky130_fd_sc_hd__o21ai_2 _33929_ (.A1(_11575_),
    .A2(_11578_),
    .B1(_11579_),
    .Y(_11580_));
 sky130_fd_sc_hd__o21ai_2 _33930_ (.A1(_11186_),
    .A2(_11180_),
    .B1(_11188_),
    .Y(_11581_));
 sky130_fd_sc_hd__buf_6 _33931_ (.A(_10598_),
    .X(_11582_));
 sky130_fd_sc_hd__buf_6 _33932_ (.A(_11179_),
    .X(_11583_));
 sky130_fd_sc_hd__a41oi_1 _33933_ (.A1(net455),
    .A2(_19674_),
    .A3(_11582_),
    .A4(_11583_),
    .B1(_11186_),
    .Y(_11584_));
 sky130_fd_sc_hd__nand2_2 _33934_ (.A(_11576_),
    .B(_11577_),
    .Y(_11585_));
 sky130_fd_sc_hd__nand2_1 _33935_ (.A(_11584_),
    .B(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__nand3_4 _33936_ (.A(_11580_),
    .B(_11581_),
    .C(_11586_),
    .Y(_11587_));
 sky130_fd_sc_hd__nand3b_2 _33937_ (.A_N(_11578_),
    .B(_11579_),
    .C(_11585_),
    .Y(_11588_));
 sky130_fd_sc_hd__buf_4 _33938_ (.A(_11189_),
    .X(_11589_));
 sky130_fd_sc_hd__a21oi_2 _33939_ (.A1(_11589_),
    .A2(_11190_),
    .B1(_11183_),
    .Y(_11590_));
 sky130_fd_sc_hd__o21ai_2 _33940_ (.A1(_11575_),
    .A2(_11578_),
    .B1(_11589_),
    .Y(_11591_));
 sky130_fd_sc_hd__nand3_4 _33941_ (.A(_11588_),
    .B(_11590_),
    .C(_11591_),
    .Y(_11592_));
 sky130_fd_sc_hd__clkbuf_4 _33942_ (.A(_18467_),
    .X(_11593_));
 sky130_fd_sc_hd__buf_6 _33943_ (.A(_11593_),
    .X(_11594_));
 sky130_fd_sc_hd__a22oi_4 _33944_ (.A1(_11594_),
    .A2(_19684_),
    .B1(_19680_),
    .B2(_19826_),
    .Y(_11595_));
 sky130_fd_sc_hd__buf_6 _33945_ (.A(_11593_),
    .X(_11596_));
 sky130_fd_sc_hd__buf_6 _33946_ (.A(_10613_),
    .X(_11597_));
 sky130_fd_sc_hd__and4_4 _33947_ (.A(_11596_),
    .B(_05162_),
    .C(_05164_),
    .D(_11597_),
    .X(_11598_));
 sky130_fd_sc_hd__nand2_2 _33948_ (.A(_19677_),
    .B(_19830_),
    .Y(_11599_));
 sky130_fd_sc_hd__o21a_2 _33949_ (.A1(_11595_),
    .A2(_11598_),
    .B1(_11599_),
    .X(_11600_));
 sky130_fd_sc_hd__nor3_4 _33950_ (.A(_11599_),
    .B(_11595_),
    .C(_11598_),
    .Y(_11601_));
 sky130_fd_sc_hd__o2bb2ai_4 _33951_ (.A1_N(_11587_),
    .A2_N(_11592_),
    .B1(_11600_),
    .B2(_11601_),
    .Y(_11602_));
 sky130_fd_sc_hd__nor2_4 _33952_ (.A(_11601_),
    .B(_11600_),
    .Y(_11603_));
 sky130_fd_sc_hd__nand3_4 _33953_ (.A(_11603_),
    .B(_11592_),
    .C(_11587_),
    .Y(_11604_));
 sky130_fd_sc_hd__nand2_1 _33954_ (.A(_11602_),
    .B(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__a21oi_4 _33955_ (.A1(_11187_),
    .A2(_11191_),
    .B1(_11196_),
    .Y(_11606_));
 sky130_fd_sc_hd__o21a_1 _33956_ (.A1(_11213_),
    .A2(_11606_),
    .B1(_11197_),
    .X(_11607_));
 sky130_fd_sc_hd__nand2_2 _33957_ (.A(_11605_),
    .B(_11607_),
    .Y(_11608_));
 sky130_fd_sc_hd__o21ai_4 _33958_ (.A1(_11213_),
    .A2(_11606_),
    .B1(_11197_),
    .Y(_11609_));
 sky130_fd_sc_hd__nand3_4 _33959_ (.A(_11609_),
    .B(_11604_),
    .C(_11602_),
    .Y(_11610_));
 sky130_fd_sc_hd__a21o_2 _33960_ (.A1(_11204_),
    .A2(_11207_),
    .B1(_11203_),
    .X(_11611_));
 sky130_fd_sc_hd__a21oi_4 _33961_ (.A1(_11608_),
    .A2(_11610_),
    .B1(_11611_),
    .Y(_11612_));
 sky130_fd_sc_hd__a21oi_4 _33962_ (.A1(_11602_),
    .A2(_11604_),
    .B1(_11609_),
    .Y(_11613_));
 sky130_fd_sc_hd__nand2_2 _33963_ (.A(_11610_),
    .B(_11611_),
    .Y(_11614_));
 sky130_fd_sc_hd__nor2_4 _33964_ (.A(_11613_),
    .B(_11614_),
    .Y(_11615_));
 sky130_fd_sc_hd__nor2_4 _33965_ (.A(_11612_),
    .B(_11615_),
    .Y(_11616_));
 sky130_fd_sc_hd__nand2_1 _33966_ (.A(_11573_),
    .B(_11616_),
    .Y(_11617_));
 sky130_fd_sc_hd__a21oi_4 _33967_ (.A1(_11028_),
    .A2(_11029_),
    .B1(_11027_),
    .Y(_11618_));
 sky130_fd_sc_hd__o21bai_2 _33968_ (.A1(_11613_),
    .A2(_11614_),
    .B1_N(_11612_),
    .Y(_11619_));
 sky130_fd_sc_hd__nand3_4 _33969_ (.A(_11619_),
    .B(_11566_),
    .C(_11572_),
    .Y(_11620_));
 sky130_fd_sc_hd__nand3_4 _33970_ (.A(_11617_),
    .B(_11618_),
    .C(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__nand3_2 _33971_ (.A(_11616_),
    .B(_11566_),
    .C(_11572_),
    .Y(_11622_));
 sky130_fd_sc_hd__o2bb2ai_2 _33972_ (.A1_N(_11572_),
    .A2_N(_11566_),
    .B1(_11612_),
    .B2(_11615_),
    .Y(_11623_));
 sky130_fd_sc_hd__o211ai_4 _33973_ (.A1(_11027_),
    .A2(_11167_),
    .B1(_11622_),
    .C1(_11623_),
    .Y(_11624_));
 sky130_fd_sc_hd__nand2_1 _33974_ (.A(_11621_),
    .B(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__nand2_2 _33975_ (.A(_11263_),
    .B(_11262_),
    .Y(_11626_));
 sky130_vsdinv _33976_ (.A(_11626_),
    .Y(_11627_));
 sky130_fd_sc_hd__nand2_2 _33977_ (.A(_11625_),
    .B(_11627_),
    .Y(_11628_));
 sky130_vsdinv _33978_ (.A(_11628_),
    .Y(_11629_));
 sky130_fd_sc_hd__nand3_4 _33979_ (.A(_11621_),
    .B(_11624_),
    .C(_11626_),
    .Y(_11630_));
 sky130_vsdinv _33980_ (.A(_11630_),
    .Y(_11631_));
 sky130_fd_sc_hd__o2bb2ai_4 _33981_ (.A1_N(_11523_),
    .A2_N(_11532_),
    .B1(_11629_),
    .B2(_11631_),
    .Y(_11632_));
 sky130_fd_sc_hd__nand2_4 _33982_ (.A(_11628_),
    .B(_11630_),
    .Y(_11633_));
 sky130_fd_sc_hd__nand3b_4 _33983_ (.A_N(_11633_),
    .B(_11532_),
    .C(_11523_),
    .Y(_11634_));
 sky130_fd_sc_hd__a21oi_4 _33984_ (.A1(_11160_),
    .A2(_11169_),
    .B1(_10955_),
    .Y(_11635_));
 sky130_fd_sc_hd__o21ai_4 _33985_ (.A1(_11278_),
    .A2(_11635_),
    .B1(_11170_),
    .Y(_11636_));
 sky130_fd_sc_hd__a21oi_4 _33986_ (.A1(_11632_),
    .A2(_11634_),
    .B1(_11636_),
    .Y(_11637_));
 sky130_fd_sc_hd__nand2_1 _33987_ (.A(_11519_),
    .B(_11522_),
    .Y(_11638_));
 sky130_fd_sc_hd__a21oi_4 _33988_ (.A1(_11638_),
    .A2(_11526_),
    .B1(_11633_),
    .Y(_11639_));
 sky130_fd_sc_hd__nand3_2 _33989_ (.A(_11176_),
    .B(_11274_),
    .C(_11271_),
    .Y(_11640_));
 sky130_fd_sc_hd__a21boi_1 _33990_ (.A1(_11532_),
    .A2(_11523_),
    .B1_N(_11633_),
    .Y(_11641_));
 sky130_fd_sc_hd__a221oi_2 _33991_ (.A1(_11639_),
    .A2(_11523_),
    .B1(_11640_),
    .B2(_11170_),
    .C1(_11641_),
    .Y(_11642_));
 sky130_fd_sc_hd__nand2_1 _33992_ (.A(_11272_),
    .B(_11270_),
    .Y(_11643_));
 sky130_vsdinv _33993_ (.A(_11223_),
    .Y(_11644_));
 sky130_fd_sc_hd__nand2_2 _33994_ (.A(_11644_),
    .B(_11220_),
    .Y(_11645_));
 sky130_fd_sc_hd__and3_2 _33995_ (.A(_11643_),
    .B(_11273_),
    .C(_11645_),
    .X(_11646_));
 sky130_fd_sc_hd__nand2_1 _33996_ (.A(_11643_),
    .B(_11273_),
    .Y(_11647_));
 sky130_fd_sc_hd__and3_2 _33997_ (.A(_11647_),
    .B(_11220_),
    .C(_11644_),
    .X(_11648_));
 sky130_fd_sc_hd__nor2_8 _33998_ (.A(_11646_),
    .B(_11648_),
    .Y(_11649_));
 sky130_fd_sc_hd__o21ai_4 _33999_ (.A1(_11637_),
    .A2(_11642_),
    .B1(_11649_),
    .Y(_11650_));
 sky130_fd_sc_hd__nand2_1 _34000_ (.A(_11280_),
    .B(_11298_),
    .Y(_11651_));
 sky130_fd_sc_hd__nand2_2 _34001_ (.A(_11651_),
    .B(_11285_),
    .Y(_11652_));
 sky130_fd_sc_hd__nand2_1 _34002_ (.A(_11632_),
    .B(_11634_),
    .Y(_11653_));
 sky130_fd_sc_hd__o21a_1 _34003_ (.A1(_11278_),
    .A2(_11635_),
    .B1(_11170_),
    .X(_11654_));
 sky130_fd_sc_hd__nand2_4 _34004_ (.A(_11653_),
    .B(_11654_),
    .Y(_11655_));
 sky130_fd_sc_hd__nand3_4 _34005_ (.A(_11636_),
    .B(_11634_),
    .C(_11632_),
    .Y(_11656_));
 sky130_fd_sc_hd__nor2_2 _34006_ (.A(_11645_),
    .B(_11647_),
    .Y(_11657_));
 sky130_fd_sc_hd__nand2_1 _34007_ (.A(_11647_),
    .B(_11645_),
    .Y(_11658_));
 sky130_vsdinv _34008_ (.A(_11658_),
    .Y(_11659_));
 sky130_fd_sc_hd__nor2_4 _34009_ (.A(_11657_),
    .B(_11659_),
    .Y(_11660_));
 sky130_fd_sc_hd__nand3_4 _34010_ (.A(_11655_),
    .B(_11656_),
    .C(_11660_),
    .Y(_11661_));
 sky130_fd_sc_hd__nand3_4 _34011_ (.A(_11650_),
    .B(_11652_),
    .C(_11661_),
    .Y(_11662_));
 sky130_fd_sc_hd__o22ai_4 _34012_ (.A1(_11646_),
    .A2(_11648_),
    .B1(_11637_),
    .B2(_11642_),
    .Y(_11663_));
 sky130_fd_sc_hd__a22oi_4 _34013_ (.A1(_11283_),
    .A2(_10903_),
    .B1(_11177_),
    .B2(_11278_),
    .Y(_11664_));
 sky130_fd_sc_hd__a22oi_4 _34014_ (.A1(_11664_),
    .A2(_11282_),
    .B1(_11280_),
    .B2(_11298_),
    .Y(_11665_));
 sky130_fd_sc_hd__nand3_4 _34015_ (.A(_11655_),
    .B(_11656_),
    .C(_11649_),
    .Y(_11666_));
 sky130_fd_sc_hd__nand3_4 _34016_ (.A(_11663_),
    .B(_11665_),
    .C(_11666_),
    .Y(_11667_));
 sky130_fd_sc_hd__nand2_1 _34017_ (.A(_11662_),
    .B(_11667_),
    .Y(_11668_));
 sky130_vsdinv _34018_ (.A(_11288_),
    .Y(_11669_));
 sky130_fd_sc_hd__a21oi_4 _34019_ (.A1(_11287_),
    .A2(_11294_),
    .B1(_11669_),
    .Y(_11670_));
 sky130_fd_sc_hd__nand2_2 _34020_ (.A(_11668_),
    .B(_11670_),
    .Y(_11671_));
 sky130_vsdinv _34021_ (.A(_11670_),
    .Y(_11672_));
 sky130_fd_sc_hd__nand3_4 _34022_ (.A(_11662_),
    .B(_11667_),
    .C(_11672_),
    .Y(_11673_));
 sky130_fd_sc_hd__nand2_2 _34023_ (.A(_11671_),
    .B(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__nand2_1 _34024_ (.A(_11301_),
    .B(_10935_),
    .Y(_11675_));
 sky130_fd_sc_hd__and2_2 _34025_ (.A(_11675_),
    .B(_11305_),
    .X(_11676_));
 sky130_fd_sc_hd__nand2_8 _34026_ (.A(_11674_),
    .B(_11676_),
    .Y(_11677_));
 sky130_fd_sc_hd__nand2_1 _34027_ (.A(_11675_),
    .B(_11305_),
    .Y(_11678_));
 sky130_fd_sc_hd__nand3_4 _34028_ (.A(_11671_),
    .B(_11678_),
    .C(_11673_),
    .Y(_11679_));
 sky130_fd_sc_hd__nand2_4 _34029_ (.A(_11677_),
    .B(_11679_),
    .Y(_11680_));
 sky130_vsdinv _34030_ (.A(_11310_),
    .Y(_11681_));
 sky130_fd_sc_hd__a21oi_4 _34031_ (.A1(net409),
    .A2(_11309_),
    .B1(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__xor2_4 _34032_ (.A(_11680_),
    .B(_11682_),
    .X(_02652_));
 sky130_fd_sc_hd__a21oi_4 _34033_ (.A1(_11655_),
    .A2(_11660_),
    .B1(_11642_),
    .Y(_11683_));
 sky130_vsdinv _34034_ (.A(_11615_),
    .Y(_11684_));
 sky130_fd_sc_hd__nand2_2 _34035_ (.A(_11684_),
    .B(_11610_),
    .Y(_11685_));
 sky130_fd_sc_hd__nand2_4 _34036_ (.A(_11630_),
    .B(_11624_),
    .Y(_11686_));
 sky130_vsdinv _34037_ (.A(_11686_),
    .Y(_11687_));
 sky130_fd_sc_hd__nor2_4 _34038_ (.A(_11685_),
    .B(_11687_),
    .Y(_11688_));
 sky130_vsdinv _34039_ (.A(_11685_),
    .Y(_11689_));
 sky130_fd_sc_hd__nor2_4 _34040_ (.A(_11689_),
    .B(_11686_),
    .Y(_11690_));
 sky130_fd_sc_hd__o21a_2 _34041_ (.A1(_11499_),
    .A2(_11469_),
    .B1(_11503_),
    .X(_11691_));
 sky130_fd_sc_hd__nand2_1 _34042_ (.A(_11460_),
    .B(_11465_),
    .Y(_11692_));
 sky130_fd_sc_hd__nand2_2 _34043_ (.A(_11692_),
    .B(_11464_),
    .Y(_11693_));
 sky130_fd_sc_hd__buf_8 _34044_ (.A(_10959_),
    .X(_11694_));
 sky130_fd_sc_hd__buf_6 _34045_ (.A(_07923_),
    .X(_11695_));
 sky130_fd_sc_hd__nand2_4 _34046_ (.A(_11695_),
    .B(_07056_),
    .Y(_11696_));
 sky130_fd_sc_hd__a21o_1 _34047_ (.A1(_10999_),
    .A2(_10733_),
    .B1(_11696_),
    .X(_11697_));
 sky130_fd_sc_hd__nand2_2 _34048_ (.A(_08623_),
    .B(_09607_),
    .Y(_11698_));
 sky130_fd_sc_hd__a21o_1 _34049_ (.A1(_10998_),
    .A2(_07344_),
    .B1(_11698_),
    .X(_11699_));
 sky130_fd_sc_hd__o211ai_4 _34050_ (.A1(net444),
    .A2(_11694_),
    .B1(_11697_),
    .C1(_11699_),
    .Y(_11700_));
 sky130_fd_sc_hd__nand3_2 _34051_ (.A(_19632_),
    .B(_19636_),
    .C(_19878_),
    .Y(_11701_));
 sky130_fd_sc_hd__nand2_1 _34052_ (.A(_11696_),
    .B(_11698_),
    .Y(_11702_));
 sky130_fd_sc_hd__o2111ai_4 _34053_ (.A1(_10724_),
    .A2(_11701_),
    .B1(net458),
    .C1(_10957_),
    .D1(_11702_),
    .Y(_11703_));
 sky130_fd_sc_hd__nand2_1 _34054_ (.A(_11700_),
    .B(_11703_),
    .Y(_11704_));
 sky130_fd_sc_hd__o21ai_2 _34055_ (.A1(_11419_),
    .A2(_11420_),
    .B1(_11422_),
    .Y(_11705_));
 sky130_fd_sc_hd__nand2_1 _34056_ (.A(_11419_),
    .B(_11420_),
    .Y(_11706_));
 sky130_fd_sc_hd__nand2_4 _34057_ (.A(_11705_),
    .B(_11706_),
    .Y(_11707_));
 sky130_fd_sc_hd__nand2_2 _34058_ (.A(_11704_),
    .B(_11707_),
    .Y(_11708_));
 sky130_fd_sc_hd__nand3b_4 _34059_ (.A_N(_11707_),
    .B(_11700_),
    .C(_11703_),
    .Y(_11709_));
 sky130_fd_sc_hd__nand2_1 _34060_ (.A(_11708_),
    .B(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__a21oi_4 _34061_ (.A1(_11452_),
    .A2(_11458_),
    .B1(_11451_),
    .Y(_11711_));
 sky130_vsdinv _34062_ (.A(_11711_),
    .Y(_11712_));
 sky130_fd_sc_hd__nand2_1 _34063_ (.A(_11710_),
    .B(_11712_),
    .Y(_11713_));
 sky130_fd_sc_hd__nand3_2 _34064_ (.A(_11708_),
    .B(_11709_),
    .C(_11711_),
    .Y(_11714_));
 sky130_fd_sc_hd__nand3b_4 _34065_ (.A_N(_11693_),
    .B(_11713_),
    .C(_11714_),
    .Y(_11715_));
 sky130_fd_sc_hd__nand2_1 _34066_ (.A(_11710_),
    .B(_11711_),
    .Y(_11716_));
 sky130_fd_sc_hd__nand3_2 _34067_ (.A(_11708_),
    .B(_11709_),
    .C(_11712_),
    .Y(_11717_));
 sky130_fd_sc_hd__nand3_4 _34068_ (.A(_11716_),
    .B(_11717_),
    .C(_11693_),
    .Y(_11718_));
 sky130_fd_sc_hd__and4_4 _34069_ (.A(_06606_),
    .B(_06907_),
    .C(_09772_),
    .D(_07705_),
    .X(_11719_));
 sky130_fd_sc_hd__a22o_2 _34070_ (.A1(_06342_),
    .A2(_10149_),
    .B1(_06343_),
    .B2(_19866_),
    .X(_11720_));
 sky130_fd_sc_hd__clkbuf_8 _34071_ (.A(_06030_),
    .X(_11721_));
 sky130_fd_sc_hd__nor2_8 _34072_ (.A(_11721_),
    .B(net439),
    .Y(_11722_));
 sky130_fd_sc_hd__nand3b_4 _34073_ (.A_N(_11719_),
    .B(_11720_),
    .C(_11722_),
    .Y(_11723_));
 sky130_fd_sc_hd__buf_4 _34074_ (.A(_10149_),
    .X(_11724_));
 sky130_fd_sc_hd__a22oi_4 _34075_ (.A1(_19645_),
    .A2(_11724_),
    .B1(_19648_),
    .B2(_10745_),
    .Y(_11725_));
 sky130_fd_sc_hd__o21bai_4 _34076_ (.A1(_11725_),
    .A2(_11719_),
    .B1_N(_11722_),
    .Y(_11726_));
 sky130_fd_sc_hd__a21o_4 _34077_ (.A1(_11474_),
    .A2(_11480_),
    .B1(_11479_),
    .X(_11727_));
 sky130_fd_sc_hd__a21o_2 _34078_ (.A1(_11723_),
    .A2(_11726_),
    .B1(_11727_),
    .X(_11728_));
 sky130_fd_sc_hd__nand3_4 _34079_ (.A(_11727_),
    .B(_11723_),
    .C(_11726_),
    .Y(_11729_));
 sky130_fd_sc_hd__nand2_1 _34080_ (.A(_11728_),
    .B(_11729_),
    .Y(_11730_));
 sky130_fd_sc_hd__nand2_1 _34081_ (.A(_06838_),
    .B(_09082_),
    .Y(_11731_));
 sky130_fd_sc_hd__nand2_1 _34082_ (.A(_06327_),
    .B(_11232_),
    .Y(_11732_));
 sky130_fd_sc_hd__a22o_1 _34083_ (.A1(_10737_),
    .A2(_19859_),
    .B1(_06336_),
    .B2(_09365_),
    .X(_11733_));
 sky130_fd_sc_hd__o21ai_1 _34084_ (.A1(_11731_),
    .A2(_11732_),
    .B1(_11733_),
    .Y(_11734_));
 sky130_fd_sc_hd__nand2_1 _34085_ (.A(_05732_),
    .B(_09823_),
    .Y(_11735_));
 sky130_fd_sc_hd__nand2_1 _34086_ (.A(_11734_),
    .B(_11735_),
    .Y(_11736_));
 sky130_fd_sc_hd__nor2_2 _34087_ (.A(_11731_),
    .B(_11732_),
    .Y(_11737_));
 sky130_vsdinv _34088_ (.A(_11735_),
    .Y(_11738_));
 sky130_fd_sc_hd__nand3b_2 _34089_ (.A_N(_11737_),
    .B(_11738_),
    .C(_11733_),
    .Y(_11739_));
 sky130_fd_sc_hd__nand2_4 _34090_ (.A(_11736_),
    .B(_11739_),
    .Y(_11740_));
 sky130_vsdinv _34091_ (.A(_11740_),
    .Y(_11741_));
 sky130_fd_sc_hd__nand2_1 _34092_ (.A(_11730_),
    .B(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__nand3_2 _34093_ (.A(_11728_),
    .B(_11729_),
    .C(_11740_),
    .Y(_11743_));
 sky130_fd_sc_hd__nand2_2 _34094_ (.A(_11742_),
    .B(_11743_),
    .Y(_11744_));
 sky130_fd_sc_hd__a21o_1 _34095_ (.A1(_11715_),
    .A2(_11718_),
    .B1(_11744_),
    .X(_11745_));
 sky130_fd_sc_hd__a21o_1 _34096_ (.A1(_11430_),
    .A2(_11431_),
    .B1(_11429_),
    .X(_11746_));
 sky130_fd_sc_hd__nand3_4 _34097_ (.A(_11715_),
    .B(_11744_),
    .C(_11718_),
    .Y(_11747_));
 sky130_fd_sc_hd__nand3_4 _34098_ (.A(_11745_),
    .B(_11746_),
    .C(_11747_),
    .Y(_11748_));
 sky130_fd_sc_hd__and2_1 _34099_ (.A(_11730_),
    .B(_11741_),
    .X(_11749_));
 sky130_vsdinv _34100_ (.A(_11743_),
    .Y(_11750_));
 sky130_fd_sc_hd__o2bb2ai_4 _34101_ (.A1_N(_11718_),
    .A2_N(_11715_),
    .B1(_11749_),
    .B2(_11750_),
    .Y(_11751_));
 sky130_fd_sc_hd__a21oi_4 _34102_ (.A1(_11430_),
    .A2(_11431_),
    .B1(_11429_),
    .Y(_11752_));
 sky130_fd_sc_hd__nand2_1 _34103_ (.A(_11730_),
    .B(_11740_),
    .Y(_11753_));
 sky130_fd_sc_hd__nand3_1 _34104_ (.A(_11741_),
    .B(_11728_),
    .C(_11729_),
    .Y(_11754_));
 sky130_fd_sc_hd__nand2_1 _34105_ (.A(_11753_),
    .B(_11754_),
    .Y(_11755_));
 sky130_fd_sc_hd__nand3_4 _34106_ (.A(_11715_),
    .B(_11755_),
    .C(_11718_),
    .Y(_11756_));
 sky130_fd_sc_hd__nand3_4 _34107_ (.A(_11751_),
    .B(_11752_),
    .C(_11756_),
    .Y(_11757_));
 sky130_fd_sc_hd__nand2_1 _34108_ (.A(_11748_),
    .B(_11757_),
    .Y(_11758_));
 sky130_fd_sc_hd__nor2_2 _34109_ (.A(_11691_),
    .B(_11758_),
    .Y(_11759_));
 sky130_vsdinv _34110_ (.A(_11691_),
    .Y(_11760_));
 sky130_fd_sc_hd__a21oi_4 _34111_ (.A1(_11748_),
    .A2(_11757_),
    .B1(_11760_),
    .Y(_11761_));
 sky130_fd_sc_hd__nand3_4 _34112_ (.A(_11075_),
    .B(_11078_),
    .C(_19923_),
    .Y(_11762_));
 sky130_fd_sc_hd__nand2_1 _34113_ (.A(_11078_),
    .B(_05263_),
    .Y(_11763_));
 sky130_fd_sc_hd__o21ai_4 _34114_ (.A1(_05229_),
    .A2(_18473_),
    .B1(_11763_),
    .Y(_11764_));
 sky130_fd_sc_hd__o21ai_2 _34115_ (.A1(_06020_),
    .A2(_11762_),
    .B1(_11764_),
    .Y(_11765_));
 sky130_fd_sc_hd__nand2_4 _34116_ (.A(_10827_),
    .B(_05272_),
    .Y(_11766_));
 sky130_fd_sc_hd__nand2_1 _34117_ (.A(_11765_),
    .B(_11766_),
    .Y(_11767_));
 sky130_vsdinv _34118_ (.A(_11766_),
    .Y(_11768_));
 sky130_fd_sc_hd__o211ai_4 _34119_ (.A1(_05128_),
    .A2(_11762_),
    .B1(_11768_),
    .C1(_11764_),
    .Y(_11769_));
 sky130_fd_sc_hd__o21bai_2 _34120_ (.A1(_11335_),
    .A2(_11334_),
    .B1_N(_11333_),
    .Y(_11770_));
 sky130_fd_sc_hd__nand3_4 _34121_ (.A(_11767_),
    .B(_11769_),
    .C(_11770_),
    .Y(_11771_));
 sky130_fd_sc_hd__nand2_1 _34122_ (.A(_11765_),
    .B(_11768_),
    .Y(_11772_));
 sky130_fd_sc_hd__o21ai_1 _34123_ (.A1(_05199_),
    .A2(_11332_),
    .B1(_11335_),
    .Y(_11773_));
 sky130_fd_sc_hd__nand2_2 _34124_ (.A(_11339_),
    .B(_11773_),
    .Y(_11774_));
 sky130_fd_sc_hd__o211ai_4 _34125_ (.A1(_05128_),
    .A2(_11762_),
    .B1(_11766_),
    .C1(_11764_),
    .Y(_11775_));
 sky130_fd_sc_hd__nand3_4 _34126_ (.A(_11772_),
    .B(_11774_),
    .C(_11775_),
    .Y(_11776_));
 sky130_fd_sc_hd__nand2_4 _34127_ (.A(_10835_),
    .B(_05267_),
    .Y(_11777_));
 sky130_fd_sc_hd__nand2_4 _34128_ (.A(\pcpi_mul.rs2[28] ),
    .B(_05277_),
    .Y(_11778_));
 sky130_fd_sc_hd__nor2_4 _34129_ (.A(_11777_),
    .B(_11778_),
    .Y(_11779_));
 sky130_fd_sc_hd__and2_1 _34130_ (.A(_11777_),
    .B(_11778_),
    .X(_11780_));
 sky130_fd_sc_hd__nand2_2 _34131_ (.A(\pcpi_mul.rs2[27] ),
    .B(_05769_),
    .Y(_11781_));
 sky130_vsdinv _34132_ (.A(_11781_),
    .Y(_11782_));
 sky130_fd_sc_hd__o21ai_2 _34133_ (.A1(_11779_),
    .A2(_11780_),
    .B1(_11782_),
    .Y(_11783_));
 sky130_vsdinv _34134_ (.A(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__or2_1 _34135_ (.A(_11777_),
    .B(_11778_),
    .X(_11785_));
 sky130_fd_sc_hd__nand2_4 _34136_ (.A(_11777_),
    .B(_11778_),
    .Y(_11786_));
 sky130_fd_sc_hd__nand3_4 _34137_ (.A(_11785_),
    .B(_11781_),
    .C(_11786_),
    .Y(_11787_));
 sky130_vsdinv _34138_ (.A(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__o2bb2ai_4 _34139_ (.A1_N(_11771_),
    .A2_N(_11776_),
    .B1(_11784_),
    .B2(_11788_),
    .Y(_11789_));
 sky130_fd_sc_hd__nand2_4 _34140_ (.A(_11783_),
    .B(_11787_),
    .Y(_11790_));
 sky130_fd_sc_hd__nand3b_4 _34141_ (.A_N(_11790_),
    .B(_11771_),
    .C(_11776_),
    .Y(_11791_));
 sky130_fd_sc_hd__a21boi_4 _34142_ (.A1(_11346_),
    .A2(_11362_),
    .B1_N(_11342_),
    .Y(_11792_));
 sky130_fd_sc_hd__nand3_4 _34143_ (.A(_11789_),
    .B(_11791_),
    .C(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__a21o_1 _34144_ (.A1(_11771_),
    .A2(_11776_),
    .B1(_11790_),
    .X(_11794_));
 sky130_fd_sc_hd__nand2_1 _34145_ (.A(_11346_),
    .B(_11362_),
    .Y(_11795_));
 sky130_fd_sc_hd__nand2_1 _34146_ (.A(_11795_),
    .B(_11342_),
    .Y(_11796_));
 sky130_fd_sc_hd__nand3_2 _34147_ (.A(_11771_),
    .B(_11776_),
    .C(_11790_),
    .Y(_11797_));
 sky130_fd_sc_hd__nand3_4 _34148_ (.A(_11794_),
    .B(_11796_),
    .C(_11797_),
    .Y(_11798_));
 sky130_fd_sc_hd__nand2_2 _34149_ (.A(_19595_),
    .B(_05660_),
    .Y(_11799_));
 sky130_fd_sc_hd__a21o_1 _34150_ (.A1(_08946_),
    .A2(_19904_),
    .B1(_11799_),
    .X(_11800_));
 sky130_fd_sc_hd__clkbuf_4 _34151_ (.A(\pcpi_mul.rs2[24] ),
    .X(_11801_));
 sky130_fd_sc_hd__nand2_1 _34152_ (.A(_11801_),
    .B(_06260_),
    .Y(_11802_));
 sky130_fd_sc_hd__nand3_2 _34153_ (.A(_11799_),
    .B(_10261_),
    .C(_06827_),
    .Y(_11803_));
 sky130_fd_sc_hd__nand3_4 _34154_ (.A(_11800_),
    .B(_11802_),
    .C(_11803_),
    .Y(_11804_));
 sky130_fd_sc_hd__nand3_2 _34155_ (.A(_19596_),
    .B(_09227_),
    .C(_06105_),
    .Y(_11805_));
 sky130_fd_sc_hd__nand2_2 _34156_ (.A(_08945_),
    .B(_05801_),
    .Y(_11806_));
 sky130_fd_sc_hd__nand2_1 _34157_ (.A(_11799_),
    .B(_11806_),
    .Y(_11807_));
 sky130_fd_sc_hd__o2111ai_4 _34158_ (.A1(_05802_),
    .A2(_11805_),
    .B1(_11801_),
    .C1(_06260_),
    .D1(_11807_),
    .Y(_11808_));
 sky130_fd_sc_hd__nand2_1 _34159_ (.A(_11804_),
    .B(_11808_),
    .Y(_11809_));
 sky130_fd_sc_hd__a21oi_2 _34160_ (.A1(_11355_),
    .A2(_11359_),
    .B1(_11353_),
    .Y(_11810_));
 sky130_fd_sc_hd__nand2_2 _34161_ (.A(_11809_),
    .B(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__nor2_2 _34162_ (.A(_11347_),
    .B(_11349_),
    .Y(_11812_));
 sky130_fd_sc_hd__o211ai_4 _34163_ (.A1(_11353_),
    .A2(_11812_),
    .B1(_11804_),
    .C1(_11808_),
    .Y(_11813_));
 sky130_fd_sc_hd__a21oi_4 _34164_ (.A1(_11376_),
    .A2(_11377_),
    .B1(_11375_),
    .Y(_11814_));
 sky130_vsdinv _34165_ (.A(_11814_),
    .Y(_11815_));
 sky130_fd_sc_hd__a21oi_4 _34166_ (.A1(_11811_),
    .A2(_11813_),
    .B1(_11815_),
    .Y(_11816_));
 sky130_fd_sc_hd__o211a_1 _34167_ (.A1(_11353_),
    .A2(_11812_),
    .B1(_11808_),
    .C1(_11804_),
    .X(_11817_));
 sky130_fd_sc_hd__nand2_1 _34168_ (.A(_11811_),
    .B(_11815_),
    .Y(_11818_));
 sky130_fd_sc_hd__nor2_1 _34169_ (.A(_11817_),
    .B(_11818_),
    .Y(_11819_));
 sky130_fd_sc_hd__o2bb2ai_2 _34170_ (.A1_N(_11793_),
    .A2_N(_11798_),
    .B1(_11816_),
    .B2(_11819_),
    .Y(_11820_));
 sky130_fd_sc_hd__nand3_2 _34171_ (.A(_11370_),
    .B(_11395_),
    .C(_11394_),
    .Y(_11821_));
 sky130_fd_sc_hd__nand2_2 _34172_ (.A(_11821_),
    .B(_11364_),
    .Y(_11822_));
 sky130_fd_sc_hd__a21boi_4 _34173_ (.A1(_11804_),
    .A2(_11808_),
    .B1_N(_11810_),
    .Y(_11823_));
 sky130_fd_sc_hd__nor2_2 _34174_ (.A(_11814_),
    .B(_11823_),
    .Y(_11824_));
 sky130_fd_sc_hd__a21oi_4 _34175_ (.A1(_11824_),
    .A2(_11813_),
    .B1(_11816_),
    .Y(_11825_));
 sky130_fd_sc_hd__nand3_4 _34176_ (.A(_11798_),
    .B(_11825_),
    .C(_11793_),
    .Y(_11826_));
 sky130_fd_sc_hd__nand3_4 _34177_ (.A(_11820_),
    .B(_11822_),
    .C(_11826_),
    .Y(_11827_));
 sky130_fd_sc_hd__nand2_1 _34178_ (.A(_11798_),
    .B(_11793_),
    .Y(_11828_));
 sky130_fd_sc_hd__nand2_1 _34179_ (.A(_11828_),
    .B(_11825_),
    .Y(_11829_));
 sky130_fd_sc_hd__a21boi_2 _34180_ (.A1(_11391_),
    .A2(_11370_),
    .B1_N(_11364_),
    .Y(_11830_));
 sky130_fd_sc_hd__nand3b_4 _34181_ (.A_N(_11825_),
    .B(_11793_),
    .C(_11798_),
    .Y(_11831_));
 sky130_fd_sc_hd__nand3_4 _34182_ (.A(_11829_),
    .B(_11830_),
    .C(_11831_),
    .Y(_11832_));
 sky130_fd_sc_hd__nand3_4 _34183_ (.A(_19607_),
    .B(_07984_),
    .C(_06657_),
    .Y(_11833_));
 sky130_fd_sc_hd__nor2_8 _34184_ (.A(net443),
    .B(_11833_),
    .Y(_11834_));
 sky130_fd_sc_hd__a22o_2 _34185_ (.A1(_08908_),
    .A2(_05774_),
    .B1(_08550_),
    .B2(_05962_),
    .X(_11835_));
 sky130_fd_sc_hd__nand2_2 _34186_ (.A(_19616_),
    .B(_06779_),
    .Y(_11836_));
 sky130_vsdinv _34187_ (.A(_11836_),
    .Y(_11837_));
 sky130_fd_sc_hd__nand3b_2 _34188_ (.A_N(_11834_),
    .B(_11835_),
    .C(_11837_),
    .Y(_11838_));
 sky130_fd_sc_hd__o21bai_2 _34189_ (.A1(_11404_),
    .A2(_11407_),
    .B1_N(_11406_),
    .Y(_11839_));
 sky130_fd_sc_hd__a22oi_4 _34190_ (.A1(_08908_),
    .A2(_06649_),
    .B1(_08550_),
    .B2(_06650_),
    .Y(_11840_));
 sky130_fd_sc_hd__o21ai_2 _34191_ (.A1(_11840_),
    .A2(_11834_),
    .B1(_11836_),
    .Y(_11841_));
 sky130_fd_sc_hd__nand3_4 _34192_ (.A(_11838_),
    .B(_11839_),
    .C(_11841_),
    .Y(_11842_));
 sky130_fd_sc_hd__o21ai_2 _34193_ (.A1(_11840_),
    .A2(_11834_),
    .B1(_11837_),
    .Y(_11843_));
 sky130_fd_sc_hd__a21oi_2 _34194_ (.A1(_11411_),
    .A2(_11410_),
    .B1(_11406_),
    .Y(_11844_));
 sky130_fd_sc_hd__o211ai_2 _34195_ (.A1(_06471_),
    .A2(_11833_),
    .B1(_11836_),
    .C1(_11835_),
    .Y(_11845_));
 sky130_fd_sc_hd__nand3_4 _34196_ (.A(_11843_),
    .B(_11844_),
    .C(_11845_),
    .Y(_11846_));
 sky130_fd_sc_hd__buf_6 _34197_ (.A(_07978_),
    .X(_11847_));
 sky130_fd_sc_hd__buf_6 _34198_ (.A(_07330_),
    .X(_11848_));
 sky130_fd_sc_hd__clkbuf_8 _34199_ (.A(_08172_),
    .X(_11849_));
 sky130_fd_sc_hd__a22oi_4 _34200_ (.A1(_11847_),
    .A2(_11848_),
    .B1(_11849_),
    .B2(_07060_),
    .Y(_11850_));
 sky130_fd_sc_hd__and4_1 _34201_ (.A(_07484_),
    .B(_07825_),
    .C(_07323_),
    .D(_07064_),
    .X(_11851_));
 sky130_fd_sc_hd__nand2_2 _34202_ (.A(_10364_),
    .B(_06799_),
    .Y(_11852_));
 sky130_vsdinv _34203_ (.A(_11852_),
    .Y(_11853_));
 sky130_fd_sc_hd__o21ai_2 _34204_ (.A1(_11850_),
    .A2(_11851_),
    .B1(_11853_),
    .Y(_11854_));
 sky130_fd_sc_hd__nand2_1 _34205_ (.A(_07484_),
    .B(_07327_),
    .Y(_11855_));
 sky130_fd_sc_hd__nand3b_4 _34206_ (.A_N(_11855_),
    .B(_19626_),
    .C(_19885_),
    .Y(_11856_));
 sky130_fd_sc_hd__a22o_1 _34207_ (.A1(_19622_),
    .A2(_06640_),
    .B1(_08565_),
    .B2(_06635_),
    .X(_11857_));
 sky130_fd_sc_hd__nand3_2 _34208_ (.A(_11856_),
    .B(_11852_),
    .C(_11857_),
    .Y(_11858_));
 sky130_fd_sc_hd__nand2_4 _34209_ (.A(_11854_),
    .B(_11858_),
    .Y(_11859_));
 sky130_fd_sc_hd__a21o_2 _34210_ (.A1(_11842_),
    .A2(_11846_),
    .B1(_11859_),
    .X(_11860_));
 sky130_fd_sc_hd__nand3_4 _34211_ (.A(_11842_),
    .B(_11846_),
    .C(_11859_),
    .Y(_11861_));
 sky130_fd_sc_hd__nand2_1 _34212_ (.A(_11860_),
    .B(_11861_),
    .Y(_11862_));
 sky130_fd_sc_hd__o21a_1 _34213_ (.A1(_11372_),
    .A2(_11384_),
    .B1(_11386_),
    .X(_11863_));
 sky130_fd_sc_hd__nand2_2 _34214_ (.A(_11862_),
    .B(_11863_),
    .Y(_11864_));
 sky130_fd_sc_hd__o21ai_4 _34215_ (.A1(_11372_),
    .A2(_11384_),
    .B1(_11386_),
    .Y(_11865_));
 sky130_fd_sc_hd__nand3_4 _34216_ (.A(_11865_),
    .B(_11860_),
    .C(_11861_),
    .Y(_11866_));
 sky130_fd_sc_hd__and2_1 _34217_ (.A(_11428_),
    .B(_11413_),
    .X(_11867_));
 sky130_fd_sc_hd__buf_2 _34218_ (.A(_11867_),
    .X(_11868_));
 sky130_vsdinv _34219_ (.A(_11868_),
    .Y(_11869_));
 sky130_fd_sc_hd__a21oi_2 _34220_ (.A1(_11864_),
    .A2(_11866_),
    .B1(_11869_),
    .Y(_11870_));
 sky130_fd_sc_hd__and3_2 _34221_ (.A(_11865_),
    .B(_11860_),
    .C(_11861_),
    .X(_11871_));
 sky130_fd_sc_hd__nand2_1 _34222_ (.A(_11869_),
    .B(_11864_),
    .Y(_11872_));
 sky130_fd_sc_hd__nor2_2 _34223_ (.A(_11871_),
    .B(_11872_),
    .Y(_11873_));
 sky130_fd_sc_hd__o2bb2ai_4 _34224_ (.A1_N(_11827_),
    .A2_N(_11832_),
    .B1(_11870_),
    .B2(_11873_),
    .Y(_11874_));
 sky130_fd_sc_hd__a21oi_4 _34225_ (.A1(_11860_),
    .A2(_11861_),
    .B1(_11865_),
    .Y(_11875_));
 sky130_fd_sc_hd__o21ai_2 _34226_ (.A1(_11875_),
    .A2(_11871_),
    .B1(_11869_),
    .Y(_11876_));
 sky130_fd_sc_hd__nand3_2 _34227_ (.A(_11864_),
    .B(_11868_),
    .C(_11866_),
    .Y(_11877_));
 sky130_fd_sc_hd__nand2_4 _34228_ (.A(_11876_),
    .B(_11877_),
    .Y(_11878_));
 sky130_fd_sc_hd__nand3_4 _34229_ (.A(_11878_),
    .B(_11827_),
    .C(_11832_),
    .Y(_11879_));
 sky130_fd_sc_hd__a21oi_2 _34230_ (.A1(_11399_),
    .A2(_11401_),
    .B1(_11400_),
    .Y(_11880_));
 sky130_fd_sc_hd__o21ai_4 _34231_ (.A1(_11435_),
    .A2(_11880_),
    .B1(_11402_),
    .Y(_11881_));
 sky130_fd_sc_hd__a21oi_4 _34232_ (.A1(_11874_),
    .A2(_11879_),
    .B1(_11881_),
    .Y(_11882_));
 sky130_vsdinv _34233_ (.A(_11402_),
    .Y(_11883_));
 sky130_fd_sc_hd__nand2_1 _34234_ (.A(_11399_),
    .B(_11401_),
    .Y(_11884_));
 sky130_fd_sc_hd__a21oi_2 _34235_ (.A1(_11884_),
    .A2(_11393_),
    .B1(_11435_),
    .Y(_11885_));
 sky130_fd_sc_hd__o211a_2 _34236_ (.A1(_11883_),
    .A2(_11885_),
    .B1(_11879_),
    .C1(_11874_),
    .X(_11886_));
 sky130_fd_sc_hd__o22ai_4 _34237_ (.A1(_11759_),
    .A2(_11761_),
    .B1(_11882_),
    .B2(_11886_),
    .Y(_11887_));
 sky130_fd_sc_hd__a21oi_1 _34238_ (.A1(_11436_),
    .A2(_11443_),
    .B1(_11441_),
    .Y(_11888_));
 sky130_fd_sc_hd__o21ai_2 _34239_ (.A1(_11529_),
    .A2(_11888_),
    .B1(_11444_),
    .Y(_11889_));
 sky130_fd_sc_hd__a21oi_2 _34240_ (.A1(_11832_),
    .A2(_11827_),
    .B1(_11878_),
    .Y(_11890_));
 sky130_fd_sc_hd__o21ai_1 _34241_ (.A1(_11875_),
    .A2(_11871_),
    .B1(_11868_),
    .Y(_11891_));
 sky130_fd_sc_hd__o2111a_1 _34242_ (.A1(_11871_),
    .A2(_11872_),
    .B1(_11891_),
    .C1(_11827_),
    .D1(_11832_),
    .X(_11892_));
 sky130_fd_sc_hd__o21bai_4 _34243_ (.A1(_11890_),
    .A2(_11892_),
    .B1_N(_11881_),
    .Y(_11893_));
 sky130_fd_sc_hd__a31oi_4 _34244_ (.A1(_11751_),
    .A2(_11752_),
    .A3(_11756_),
    .B1(_11691_),
    .Y(_11894_));
 sky130_fd_sc_hd__a21oi_4 _34245_ (.A1(_11748_),
    .A2(_11894_),
    .B1(_11761_),
    .Y(_11895_));
 sky130_fd_sc_hd__nand3_4 _34246_ (.A(_11881_),
    .B(_11874_),
    .C(_11879_),
    .Y(_11896_));
 sky130_fd_sc_hd__nand3_2 _34247_ (.A(_11893_),
    .B(_11895_),
    .C(_11896_),
    .Y(_11897_));
 sky130_fd_sc_hd__nand3_4 _34248_ (.A(_11887_),
    .B(_11889_),
    .C(_11897_),
    .Y(_11898_));
 sky130_fd_sc_hd__o21ai_2 _34249_ (.A1(_11882_),
    .A2(_11886_),
    .B1(_11895_),
    .Y(_11899_));
 sky130_fd_sc_hd__a21boi_4 _34250_ (.A1(_11521_),
    .A2(_11448_),
    .B1_N(_11444_),
    .Y(_11900_));
 sky130_fd_sc_hd__nand2_1 _34251_ (.A(_11758_),
    .B(_11691_),
    .Y(_11901_));
 sky130_fd_sc_hd__nand2_1 _34252_ (.A(_11894_),
    .B(_11748_),
    .Y(_11902_));
 sky130_fd_sc_hd__nand2_2 _34253_ (.A(_11901_),
    .B(_11902_),
    .Y(_11903_));
 sky130_fd_sc_hd__nand3_4 _34254_ (.A(_11893_),
    .B(_11896_),
    .C(_11903_),
    .Y(_11904_));
 sky130_fd_sc_hd__nand3_4 _34255_ (.A(_11899_),
    .B(_11900_),
    .C(_11904_),
    .Y(_11905_));
 sky130_vsdinv _34256_ (.A(_11552_),
    .Y(_11906_));
 sky130_vsdinv _34257_ (.A(_11556_),
    .Y(_11907_));
 sky130_fd_sc_hd__and4_4 _34258_ (.A(_05841_),
    .B(_05589_),
    .C(_09817_),
    .D(_11228_),
    .X(_11908_));
 sky130_fd_sc_hd__buf_6 _34259_ (.A(_09358_),
    .X(_11909_));
 sky130_fd_sc_hd__a22o_2 _34260_ (.A1(_06493_),
    .A2(_11909_),
    .B1(_19666_),
    .B2(_19844_),
    .X(_11910_));
 sky130_fd_sc_hd__nand2_2 _34261_ (.A(_19668_),
    .B(_19839_),
    .Y(_11911_));
 sky130_vsdinv _34262_ (.A(_11911_),
    .Y(_11912_));
 sky130_fd_sc_hd__nand3b_2 _34263_ (.A_N(_11908_),
    .B(_11910_),
    .C(_11912_),
    .Y(_11913_));
 sky130_fd_sc_hd__o21bai_2 _34264_ (.A1(_11487_),
    .A2(_11484_),
    .B1_N(_11485_),
    .Y(_11914_));
 sky130_fd_sc_hd__a22oi_4 _34265_ (.A1(_06493_),
    .A2(_11909_),
    .B1(_06505_),
    .B2(_11178_),
    .Y(_11915_));
 sky130_fd_sc_hd__o21ai_2 _34266_ (.A1(_11915_),
    .A2(_11908_),
    .B1(_11911_),
    .Y(_11916_));
 sky130_fd_sc_hd__nand3_4 _34267_ (.A(_11913_),
    .B(_11914_),
    .C(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__nor2_1 _34268_ (.A(_11487_),
    .B(_11484_),
    .Y(_11918_));
 sky130_fd_sc_hd__nor2_2 _34269_ (.A(_11485_),
    .B(_11918_),
    .Y(_11919_));
 sky130_fd_sc_hd__nand3b_2 _34270_ (.A_N(_11908_),
    .B(_11910_),
    .C(_11911_),
    .Y(_11920_));
 sky130_fd_sc_hd__o21ai_2 _34271_ (.A1(_11915_),
    .A2(_11908_),
    .B1(_11912_),
    .Y(_11921_));
 sky130_fd_sc_hd__nand3_4 _34272_ (.A(_11919_),
    .B(_11920_),
    .C(_11921_),
    .Y(_11922_));
 sky130_fd_sc_hd__nor2_8 _34273_ (.A(_11541_),
    .B(_11539_),
    .Y(_11923_));
 sky130_fd_sc_hd__o2bb2ai_4 _34274_ (.A1_N(_11917_),
    .A2_N(_11922_),
    .B1(_11535_),
    .B2(_11923_),
    .Y(_11924_));
 sky130_fd_sc_hd__nor2_4 _34275_ (.A(_11535_),
    .B(_11923_),
    .Y(_11925_));
 sky130_fd_sc_hd__nand3_4 _34276_ (.A(_11922_),
    .B(_11917_),
    .C(_11925_),
    .Y(_11926_));
 sky130_fd_sc_hd__nand2_4 _34277_ (.A(_11495_),
    .B(_11482_),
    .Y(_11927_));
 sky130_fd_sc_hd__a21oi_4 _34278_ (.A1(_11924_),
    .A2(_11926_),
    .B1(_11927_),
    .Y(_11928_));
 sky130_fd_sc_hd__and3_1 _34279_ (.A(_11927_),
    .B(_11924_),
    .C(_11926_),
    .X(_11929_));
 sky130_fd_sc_hd__o22ai_4 _34280_ (.A1(_11906_),
    .A2(_11907_),
    .B1(_11928_),
    .B2(_11929_),
    .Y(_11930_));
 sky130_fd_sc_hd__nand2_1 _34281_ (.A(_11556_),
    .B(_11552_),
    .Y(_11931_));
 sky130_vsdinv _34282_ (.A(_11931_),
    .Y(_11932_));
 sky130_fd_sc_hd__nand3_4 _34283_ (.A(_11927_),
    .B(_11924_),
    .C(_11926_),
    .Y(_11933_));
 sky130_fd_sc_hd__nand3b_2 _34284_ (.A_N(_11928_),
    .B(_11932_),
    .C(_11933_),
    .Y(_11934_));
 sky130_fd_sc_hd__o21a_1 _34285_ (.A1(_11564_),
    .A2(_11558_),
    .B1(_11563_),
    .X(_11935_));
 sky130_fd_sc_hd__nand3_4 _34286_ (.A(_11930_),
    .B(_11934_),
    .C(_11935_),
    .Y(_11936_));
 sky130_fd_sc_hd__o21ai_2 _34287_ (.A1(_11928_),
    .A2(_11929_),
    .B1(_11932_),
    .Y(_11937_));
 sky130_fd_sc_hd__o21ai_2 _34288_ (.A1(_11564_),
    .A2(_11558_),
    .B1(_11563_),
    .Y(_11938_));
 sky130_fd_sc_hd__nand3b_2 _34289_ (.A_N(_11928_),
    .B(_11931_),
    .C(_11933_),
    .Y(_11939_));
 sky130_fd_sc_hd__nand3_4 _34290_ (.A(_11937_),
    .B(_11938_),
    .C(_11939_),
    .Y(_11940_));
 sky130_fd_sc_hd__nand2_2 _34291_ (.A(_05791_),
    .B(_10487_),
    .Y(_11941_));
 sky130_fd_sc_hd__nand2_2 _34292_ (.A(_05792_),
    .B(_11202_),
    .Y(_11942_));
 sky130_fd_sc_hd__or2_4 _34293_ (.A(_11941_),
    .B(_11942_),
    .X(_11943_));
 sky130_fd_sc_hd__nand2_4 _34294_ (.A(_11941_),
    .B(_11942_),
    .Y(_11944_));
 sky130_fd_sc_hd__a21o_1 _34295_ (.A1(_11943_),
    .A2(_11944_),
    .B1(_11579_),
    .X(_11945_));
 sky130_fd_sc_hd__a21oi_4 _34296_ (.A1(_11589_),
    .A2(_11585_),
    .B1(_11578_),
    .Y(_11946_));
 sky130_fd_sc_hd__nand3_2 _34297_ (.A(_11943_),
    .B(_11579_),
    .C(_11944_),
    .Y(_11947_));
 sky130_fd_sc_hd__nand3_4 _34298_ (.A(_11945_),
    .B(_11946_),
    .C(_11947_),
    .Y(_11948_));
 sky130_fd_sc_hd__o2bb2ai_2 _34299_ (.A1_N(_11944_),
    .A2_N(_11943_),
    .B1(_18469_),
    .B2(net474),
    .Y(_11949_));
 sky130_vsdinv _34300_ (.A(_11946_),
    .Y(_11950_));
 sky130_fd_sc_hd__nand3_4 _34301_ (.A(_11943_),
    .B(_11589_),
    .C(_11944_),
    .Y(_11951_));
 sky130_fd_sc_hd__nand3_4 _34302_ (.A(_11949_),
    .B(_11950_),
    .C(_11951_),
    .Y(_11952_));
 sky130_fd_sc_hd__nand2_1 _34303_ (.A(_11948_),
    .B(_11952_),
    .Y(_11953_));
 sky130_fd_sc_hd__nand2_1 _34304_ (.A(_19677_),
    .B(_19827_),
    .Y(_11954_));
 sky130_fd_sc_hd__o21ai_1 _34305_ (.A1(_19680_),
    .A2(_19684_),
    .B1(_11594_),
    .Y(_11955_));
 sky130_fd_sc_hd__nand3_4 _34306_ (.A(_18467_),
    .B(_19678_),
    .C(_19681_),
    .Y(_11956_));
 sky130_vsdinv _34307_ (.A(_11956_),
    .Y(_11957_));
 sky130_fd_sc_hd__nor2_1 _34308_ (.A(_11955_),
    .B(_11957_),
    .Y(_11958_));
 sky130_fd_sc_hd__nor2_1 _34309_ (.A(_11954_),
    .B(_11958_),
    .Y(_11959_));
 sky130_fd_sc_hd__nand2_1 _34310_ (.A(_11958_),
    .B(_11954_),
    .Y(_11960_));
 sky130_fd_sc_hd__and2b_1 _34311_ (.A_N(_11959_),
    .B(_11960_),
    .X(_11961_));
 sky130_fd_sc_hd__nand2_4 _34312_ (.A(_11953_),
    .B(_11961_),
    .Y(_11962_));
 sky130_fd_sc_hd__or2b_2 _34313_ (.A(_11959_),
    .B_N(_11960_),
    .X(_11963_));
 sky130_fd_sc_hd__nand3_4 _34314_ (.A(_11963_),
    .B(_11948_),
    .C(_11952_),
    .Y(_11964_));
 sky130_fd_sc_hd__nand2_1 _34315_ (.A(_11962_),
    .B(_11964_),
    .Y(_11965_));
 sky130_fd_sc_hd__a21boi_1 _34316_ (.A1(_11603_),
    .A2(_11592_),
    .B1_N(_11587_),
    .Y(_11966_));
 sky130_fd_sc_hd__nand2_1 _34317_ (.A(_11965_),
    .B(_11966_),
    .Y(_11967_));
 sky130_fd_sc_hd__a21bo_2 _34318_ (.A1(_11603_),
    .A2(_11592_),
    .B1_N(_11587_),
    .X(_11968_));
 sky130_fd_sc_hd__nand3_4 _34319_ (.A(_11962_),
    .B(_11968_),
    .C(_11964_),
    .Y(_11969_));
 sky130_fd_sc_hd__nor2_4 _34320_ (.A(_11598_),
    .B(_11601_),
    .Y(_11970_));
 sky130_vsdinv _34321_ (.A(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__a21oi_1 _34322_ (.A1(_11967_),
    .A2(_11969_),
    .B1(_11971_),
    .Y(_11972_));
 sky130_fd_sc_hd__and3_1 _34323_ (.A(_11967_),
    .B(_11969_),
    .C(_11971_),
    .X(_11973_));
 sky130_fd_sc_hd__o2bb2ai_2 _34324_ (.A1_N(_11936_),
    .A2_N(_11940_),
    .B1(_11972_),
    .B2(_11973_),
    .Y(_11974_));
 sky130_fd_sc_hd__a21oi_4 _34325_ (.A1(_11962_),
    .A2(_11964_),
    .B1(_11968_),
    .Y(_11975_));
 sky130_fd_sc_hd__and3_1 _34326_ (.A(_11949_),
    .B(_11950_),
    .C(_11951_),
    .X(_11976_));
 sky130_fd_sc_hd__nand2_1 _34327_ (.A(_11963_),
    .B(_11948_),
    .Y(_11977_));
 sky130_fd_sc_hd__o211a_2 _34328_ (.A1(_11976_),
    .A2(_11977_),
    .B1(_11968_),
    .C1(_11962_),
    .X(_11978_));
 sky130_fd_sc_hd__o22ai_4 _34329_ (.A1(_11598_),
    .A2(_11601_),
    .B1(_11975_),
    .B2(_11978_),
    .Y(_11979_));
 sky130_fd_sc_hd__nand3_2 _34330_ (.A(_11967_),
    .B(_11969_),
    .C(_11970_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand2_4 _34331_ (.A(_11979_),
    .B(_11980_),
    .Y(_11981_));
 sky130_fd_sc_hd__nand3_4 _34332_ (.A(_11981_),
    .B(_11936_),
    .C(_11940_),
    .Y(_11982_));
 sky130_fd_sc_hd__nand2_2 _34333_ (.A(_11514_),
    .B(_11517_),
    .Y(_11983_));
 sky130_fd_sc_hd__nand2_2 _34334_ (.A(_11983_),
    .B(_11506_),
    .Y(_11984_));
 sky130_fd_sc_hd__a21o_1 _34335_ (.A1(_11974_),
    .A2(_11982_),
    .B1(_11984_),
    .X(_11985_));
 sky130_fd_sc_hd__nand2_1 _34336_ (.A(_11940_),
    .B(_11936_),
    .Y(_11986_));
 sky130_fd_sc_hd__nor2_2 _34337_ (.A(_11970_),
    .B(_11975_),
    .Y(_11987_));
 sky130_fd_sc_hd__nand2_1 _34338_ (.A(_11987_),
    .B(_11969_),
    .Y(_11988_));
 sky130_fd_sc_hd__o21ai_1 _34339_ (.A1(_11975_),
    .A2(_11978_),
    .B1(_11970_),
    .Y(_11989_));
 sky130_fd_sc_hd__nand2_2 _34340_ (.A(_11988_),
    .B(_11989_),
    .Y(_11990_));
 sky130_fd_sc_hd__a22oi_4 _34341_ (.A1(_11983_),
    .A2(_11506_),
    .B1(_11986_),
    .B2(_11990_),
    .Y(_11991_));
 sky130_fd_sc_hd__nand2_2 _34342_ (.A(_11991_),
    .B(_11982_),
    .Y(_11992_));
 sky130_vsdinv _34343_ (.A(_11572_),
    .Y(_11993_));
 sky130_fd_sc_hd__a21o_2 _34344_ (.A1(_11566_),
    .A2(_11616_),
    .B1(_11993_),
    .X(_11994_));
 sky130_fd_sc_hd__a21oi_2 _34345_ (.A1(_11985_),
    .A2(_11992_),
    .B1(_11994_),
    .Y(_11995_));
 sky130_fd_sc_hd__and3_1 _34346_ (.A(_11974_),
    .B(_11984_),
    .C(_11982_),
    .X(_11996_));
 sky130_fd_sc_hd__nand2_1 _34347_ (.A(_11985_),
    .B(_11994_),
    .Y(_11997_));
 sky130_fd_sc_hd__nor2_2 _34348_ (.A(_11996_),
    .B(_11997_),
    .Y(_11998_));
 sky130_fd_sc_hd__o2bb2ai_4 _34349_ (.A1_N(_11898_),
    .A2_N(_11905_),
    .B1(_11995_),
    .B2(_11998_),
    .Y(_11999_));
 sky130_fd_sc_hd__and2_1 _34350_ (.A(_11616_),
    .B(_11566_),
    .X(_12000_));
 sky130_fd_sc_hd__a21oi_4 _34351_ (.A1(_11974_),
    .A2(_11982_),
    .B1(_11984_),
    .Y(_12001_));
 sky130_fd_sc_hd__o22ai_4 _34352_ (.A1(_11993_),
    .A2(_12000_),
    .B1(_12001_),
    .B2(_11996_),
    .Y(_12002_));
 sky130_vsdinv _34353_ (.A(_11994_),
    .Y(_12003_));
 sky130_fd_sc_hd__nand3_2 _34354_ (.A(_11985_),
    .B(_11992_),
    .C(_12003_),
    .Y(_12004_));
 sky130_fd_sc_hd__nand2_2 _34355_ (.A(_12002_),
    .B(_12004_),
    .Y(_12005_));
 sky130_fd_sc_hd__nand3_4 _34356_ (.A(_12005_),
    .B(_11905_),
    .C(_11898_),
    .Y(_12006_));
 sky130_fd_sc_hd__a21oi_2 _34357_ (.A1(_11519_),
    .A2(_11522_),
    .B1(_11328_),
    .Y(_12007_));
 sky130_fd_sc_hd__o21ai_4 _34358_ (.A1(_11633_),
    .A2(_12007_),
    .B1(_11523_),
    .Y(_12008_));
 sky130_fd_sc_hd__a21oi_4 _34359_ (.A1(_11999_),
    .A2(_12006_),
    .B1(_12008_),
    .Y(_12009_));
 sky130_vsdinv _34360_ (.A(_11523_),
    .Y(_12010_));
 sky130_fd_sc_hd__o211a_4 _34361_ (.A1(_12010_),
    .A2(_11639_),
    .B1(_12006_),
    .C1(_11999_),
    .X(_12011_));
 sky130_fd_sc_hd__o22ai_4 _34362_ (.A1(_11688_),
    .A2(_11690_),
    .B1(_12009_),
    .B2(_12011_),
    .Y(_12012_));
 sky130_fd_sc_hd__a21oi_2 _34363_ (.A1(_11905_),
    .A2(_11898_),
    .B1(_12005_),
    .Y(_12013_));
 sky130_fd_sc_hd__a211oi_4 _34364_ (.A1(_11991_),
    .A2(_11982_),
    .B1(_11994_),
    .C1(_12001_),
    .Y(_12014_));
 sky130_fd_sc_hd__a21oi_1 _34365_ (.A1(_11985_),
    .A2(_11992_),
    .B1(_12003_),
    .Y(_12015_));
 sky130_fd_sc_hd__o211a_1 _34366_ (.A1(_12014_),
    .A2(_12015_),
    .B1(_11898_),
    .C1(_11905_),
    .X(_12016_));
 sky130_fd_sc_hd__o21bai_4 _34367_ (.A1(_12013_),
    .A2(_12016_),
    .B1_N(_12008_),
    .Y(_12017_));
 sky130_fd_sc_hd__nand3_4 _34368_ (.A(_11999_),
    .B(_12008_),
    .C(_12006_),
    .Y(_12018_));
 sky130_fd_sc_hd__nor2_4 _34369_ (.A(_11690_),
    .B(_11688_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand3_4 _34370_ (.A(_12017_),
    .B(_12018_),
    .C(_12019_),
    .Y(_12020_));
 sky130_fd_sc_hd__nand3_4 _34371_ (.A(_11683_),
    .B(_12012_),
    .C(_12020_),
    .Y(_12021_));
 sky130_fd_sc_hd__nor2_8 _34372_ (.A(_11689_),
    .B(_11687_),
    .Y(_12022_));
 sky130_fd_sc_hd__nor2_4 _34373_ (.A(_11685_),
    .B(_11686_),
    .Y(_12023_));
 sky130_fd_sc_hd__o22ai_4 _34374_ (.A1(_12022_),
    .A2(_12023_),
    .B1(_12009_),
    .B2(_12011_),
    .Y(_12024_));
 sky130_fd_sc_hd__o21ai_2 _34375_ (.A1(_11649_),
    .A2(_11637_),
    .B1(_11656_),
    .Y(_12025_));
 sky130_fd_sc_hd__nor2_4 _34376_ (.A(_12023_),
    .B(_12022_),
    .Y(_12026_));
 sky130_fd_sc_hd__nand3_4 _34377_ (.A(_12017_),
    .B(_12018_),
    .C(_12026_),
    .Y(_12027_));
 sky130_fd_sc_hd__nand3_4 _34378_ (.A(_12024_),
    .B(_12025_),
    .C(_12027_),
    .Y(_12028_));
 sky130_fd_sc_hd__a21oi_2 _34379_ (.A1(_12021_),
    .A2(_12028_),
    .B1(_11659_),
    .Y(_12029_));
 sky130_fd_sc_hd__and3_1 _34380_ (.A(_12021_),
    .B(_12028_),
    .C(_11659_),
    .X(_12030_));
 sky130_vsdinv _34381_ (.A(_11661_),
    .Y(_12031_));
 sky130_fd_sc_hd__nand2_1 _34382_ (.A(_11650_),
    .B(_11652_),
    .Y(_12032_));
 sky130_fd_sc_hd__o2bb2ai_4 _34383_ (.A1_N(_11667_),
    .A2_N(_11672_),
    .B1(_12031_),
    .B2(_12032_),
    .Y(_12033_));
 sky130_fd_sc_hd__o21bai_4 _34384_ (.A1(_12029_),
    .A2(_12030_),
    .B1_N(_12033_),
    .Y(_12034_));
 sky130_vsdinv _34385_ (.A(_12028_),
    .Y(_12035_));
 sky130_fd_sc_hd__nand2_2 _34386_ (.A(_12021_),
    .B(_11659_),
    .Y(_12036_));
 sky130_fd_sc_hd__a21o_1 _34387_ (.A1(_12021_),
    .A2(_12028_),
    .B1(_11659_),
    .X(_12037_));
 sky130_fd_sc_hd__o211ai_4 _34388_ (.A1(_12035_),
    .A2(_12036_),
    .B1(_12033_),
    .C1(_12037_),
    .Y(_12038_));
 sky130_fd_sc_hd__and2_2 _34389_ (.A(_12034_),
    .B(_12038_),
    .X(_12039_));
 sky130_fd_sc_hd__nand2_4 _34390_ (.A(_11679_),
    .B(_11310_),
    .Y(_12040_));
 sky130_fd_sc_hd__nor2_8 _34391_ (.A(_11311_),
    .B(_11680_),
    .Y(_12041_));
 sky130_fd_sc_hd__a22oi_4 _34392_ (.A1(_11677_),
    .A2(_12040_),
    .B1(net409),
    .B2(_12041_),
    .Y(_12042_));
 sky130_fd_sc_hd__xnor2_4 _34393_ (.A(_12039_),
    .B(_12042_),
    .Y(_02653_));
 sky130_fd_sc_hd__a21oi_1 _34394_ (.A1(_11862_),
    .A2(_11863_),
    .B1(_11868_),
    .Y(_12043_));
 sky130_fd_sc_hd__a22oi_4 _34395_ (.A1(_19632_),
    .A2(_07346_),
    .B1(_19636_),
    .B2(_08062_),
    .Y(_12044_));
 sky130_fd_sc_hd__nand3_4 _34396_ (.A(_06924_),
    .B(_06921_),
    .C(_09607_),
    .Y(_12045_));
 sky130_fd_sc_hd__nor2_4 _34397_ (.A(_10960_),
    .B(_12045_),
    .Y(_12046_));
 sky130_fd_sc_hd__nand2_2 _34398_ (.A(_19641_),
    .B(_10395_),
    .Y(_12047_));
 sky130_vsdinv _34399_ (.A(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__o21ai_2 _34400_ (.A1(_12044_),
    .A2(_12046_),
    .B1(_12048_),
    .Y(_12049_));
 sky130_fd_sc_hd__a21oi_2 _34401_ (.A1(_11857_),
    .A2(_11853_),
    .B1(_11851_),
    .Y(_12050_));
 sky130_fd_sc_hd__a22o_2 _34402_ (.A1(_10998_),
    .A2(_07346_),
    .B1(_10999_),
    .B2(_08062_),
    .X(_12051_));
 sky130_fd_sc_hd__o211ai_4 _34403_ (.A1(_11694_),
    .A2(_12045_),
    .B1(_12047_),
    .C1(_12051_),
    .Y(_12052_));
 sky130_fd_sc_hd__nand3_4 _34404_ (.A(_12049_),
    .B(_12050_),
    .C(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__o21ai_2 _34405_ (.A1(_12044_),
    .A2(_12046_),
    .B1(_12047_),
    .Y(_12054_));
 sky130_fd_sc_hd__o211ai_4 _34406_ (.A1(_11694_),
    .A2(_12045_),
    .B1(_12048_),
    .C1(_12051_),
    .Y(_12055_));
 sky130_fd_sc_hd__o21ai_2 _34407_ (.A1(_11852_),
    .A2(_11850_),
    .B1(_11856_),
    .Y(_12056_));
 sky130_fd_sc_hd__nand3_4 _34408_ (.A(_12054_),
    .B(_12055_),
    .C(_12056_),
    .Y(_12057_));
 sky130_fd_sc_hd__o21ai_4 _34409_ (.A1(_11696_),
    .A2(_11698_),
    .B1(_11703_),
    .Y(_12058_));
 sky130_fd_sc_hd__nand3_4 _34410_ (.A(_12053_),
    .B(_12057_),
    .C(_12058_),
    .Y(_12059_));
 sky130_fd_sc_hd__a21o_4 _34411_ (.A1(_12053_),
    .A2(_12057_),
    .B1(_12058_),
    .X(_12060_));
 sky130_fd_sc_hd__a21boi_4 _34412_ (.A1(_11700_),
    .A2(_11703_),
    .B1_N(_11707_),
    .Y(_12061_));
 sky130_fd_sc_hd__o21a_1 _34413_ (.A1(_11707_),
    .A2(_11704_),
    .B1(_11711_),
    .X(_12062_));
 sky130_fd_sc_hd__o2bb2ai_4 _34414_ (.A1_N(_12059_),
    .A2_N(_12060_),
    .B1(_12061_),
    .B2(_12062_),
    .Y(_12063_));
 sky130_fd_sc_hd__o21ai_4 _34415_ (.A1(_11711_),
    .A2(_12061_),
    .B1(_11709_),
    .Y(_12064_));
 sky130_fd_sc_hd__nand3_4 _34416_ (.A(_12064_),
    .B(_12060_),
    .C(_12059_),
    .Y(_12065_));
 sky130_fd_sc_hd__a21o_1 _34417_ (.A1(_11722_),
    .A2(_11720_),
    .B1(_11719_),
    .X(_12066_));
 sky130_fd_sc_hd__nand3_4 _34418_ (.A(_07007_),
    .B(_06906_),
    .C(_07686_),
    .Y(_12067_));
 sky130_fd_sc_hd__nor2_8 _34419_ (.A(_08042_),
    .B(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__a22o_4 _34420_ (.A1(_06414_),
    .A2(_19865_),
    .B1(_06610_),
    .B2(_08331_),
    .X(_12069_));
 sky130_fd_sc_hd__nand2_4 _34421_ (.A(_07223_),
    .B(\pcpi_mul.rs1[23] ),
    .Y(_12070_));
 sky130_vsdinv _34422_ (.A(_12070_),
    .Y(_12071_));
 sky130_fd_sc_hd__nand3b_4 _34423_ (.A_N(_12068_),
    .B(_12069_),
    .C(_12071_),
    .Y(_12072_));
 sky130_fd_sc_hd__a22oi_4 _34424_ (.A1(net445),
    .A2(_10738_),
    .B1(_06423_),
    .B2(_19863_),
    .Y(_12073_));
 sky130_fd_sc_hd__o21ai_2 _34425_ (.A1(_12073_),
    .A2(_12068_),
    .B1(_12070_),
    .Y(_12074_));
 sky130_fd_sc_hd__nand3_4 _34426_ (.A(_12066_),
    .B(_12072_),
    .C(_12074_),
    .Y(_12075_));
 sky130_fd_sc_hd__a21oi_4 _34427_ (.A1(_11722_),
    .A2(_11720_),
    .B1(_11719_),
    .Y(_12076_));
 sky130_fd_sc_hd__o21ai_4 _34428_ (.A1(_12073_),
    .A2(_12068_),
    .B1(_12071_),
    .Y(_12077_));
 sky130_fd_sc_hd__buf_6 _34429_ (.A(_08043_),
    .X(_12078_));
 sky130_fd_sc_hd__o211ai_4 _34430_ (.A1(_12078_),
    .A2(_12067_),
    .B1(_12070_),
    .C1(_12069_),
    .Y(_12079_));
 sky130_fd_sc_hd__nand2_4 _34431_ (.A(_05883_),
    .B(_10643_),
    .Y(_12080_));
 sky130_fd_sc_hd__nand2_2 _34432_ (.A(net477),
    .B(_19851_),
    .Y(_12081_));
 sky130_fd_sc_hd__nor2_4 _34433_ (.A(_12080_),
    .B(_12081_),
    .Y(_12082_));
 sky130_fd_sc_hd__nand2_4 _34434_ (.A(_06014_),
    .B(_09820_),
    .Y(_12083_));
 sky130_fd_sc_hd__a22o_1 _34435_ (.A1(_10737_),
    .A2(_11232_),
    .B1(_06336_),
    .B2(_11224_),
    .X(_12084_));
 sky130_fd_sc_hd__nand3b_4 _34436_ (.A_N(_12082_),
    .B(_12083_),
    .C(_12084_),
    .Y(_12085_));
 sky130_fd_sc_hd__a22oi_4 _34437_ (.A1(_10737_),
    .A2(_09365_),
    .B1(_06160_),
    .B2(_11224_),
    .Y(_12086_));
 sky130_vsdinv _34438_ (.A(_12083_),
    .Y(_12087_));
 sky130_fd_sc_hd__o21ai_4 _34439_ (.A1(_12086_),
    .A2(_12082_),
    .B1(_12087_),
    .Y(_12088_));
 sky130_fd_sc_hd__a32oi_4 _34440_ (.A1(_12076_),
    .A2(_12077_),
    .A3(_12079_),
    .B1(_12085_),
    .B2(_12088_),
    .Y(_12089_));
 sky130_fd_sc_hd__nand3_4 _34441_ (.A(_12076_),
    .B(_12077_),
    .C(_12079_),
    .Y(_12090_));
 sky130_fd_sc_hd__nand2_4 _34442_ (.A(_12085_),
    .B(_12088_),
    .Y(_12091_));
 sky130_fd_sc_hd__a21oi_4 _34443_ (.A1(_12075_),
    .A2(_12090_),
    .B1(_12091_),
    .Y(_12092_));
 sky130_fd_sc_hd__a21oi_4 _34444_ (.A1(_12075_),
    .A2(_12089_),
    .B1(_12092_),
    .Y(_12093_));
 sky130_fd_sc_hd__nand3_4 _34445_ (.A(_12063_),
    .B(_12065_),
    .C(_12093_),
    .Y(_12094_));
 sky130_fd_sc_hd__nand2_1 _34446_ (.A(_12089_),
    .B(_12075_),
    .Y(_12095_));
 sky130_vsdinv _34447_ (.A(_12095_),
    .Y(_12096_));
 sky130_fd_sc_hd__o2bb2ai_4 _34448_ (.A1_N(_12065_),
    .A2_N(_12063_),
    .B1(_12092_),
    .B2(_12096_),
    .Y(_12097_));
 sky130_fd_sc_hd__o211a_2 _34449_ (.A1(_11871_),
    .A2(_12043_),
    .B1(_12094_),
    .C1(_12097_),
    .X(_12098_));
 sky130_fd_sc_hd__and2_1 _34450_ (.A(_11866_),
    .B(_11868_),
    .X(_12099_));
 sky130_fd_sc_hd__a21oi_4 _34451_ (.A1(_12063_),
    .A2(_12065_),
    .B1(_12093_),
    .Y(_12100_));
 sky130_fd_sc_hd__nand2_1 _34452_ (.A(_12075_),
    .B(_12090_),
    .Y(_12101_));
 sky130_vsdinv _34453_ (.A(_12091_),
    .Y(_12102_));
 sky130_fd_sc_hd__nand2_1 _34454_ (.A(_12101_),
    .B(_12102_),
    .Y(_12103_));
 sky130_fd_sc_hd__nand2_2 _34455_ (.A(_12095_),
    .B(_12103_),
    .Y(_12104_));
 sky130_fd_sc_hd__a21oi_4 _34456_ (.A1(_12060_),
    .A2(_12059_),
    .B1(_12064_),
    .Y(_12105_));
 sky130_fd_sc_hd__nor3b_4 _34457_ (.A(_12104_),
    .B(_12105_),
    .C_N(_12065_),
    .Y(_12106_));
 sky130_fd_sc_hd__o22ai_4 _34458_ (.A1(_11875_),
    .A2(_12099_),
    .B1(_12100_),
    .B2(_12106_),
    .Y(_12107_));
 sky130_fd_sc_hd__nand2_1 _34459_ (.A(_11715_),
    .B(_11744_),
    .Y(_12108_));
 sky130_fd_sc_hd__nand2_2 _34460_ (.A(_12108_),
    .B(_11718_),
    .Y(_12109_));
 sky130_fd_sc_hd__nand2_2 _34461_ (.A(_12107_),
    .B(_12109_),
    .Y(_12110_));
 sky130_fd_sc_hd__nor2_2 _34462_ (.A(_12098_),
    .B(_12110_),
    .Y(_12111_));
 sky130_fd_sc_hd__o21ai_4 _34463_ (.A1(_11868_),
    .A2(_11875_),
    .B1(_11866_),
    .Y(_12112_));
 sky130_fd_sc_hd__nand3_4 _34464_ (.A(_12097_),
    .B(_12112_),
    .C(_12094_),
    .Y(_12113_));
 sky130_fd_sc_hd__a21oi_4 _34465_ (.A1(_12107_),
    .A2(_12113_),
    .B1(_12109_),
    .Y(_12114_));
 sky130_fd_sc_hd__nand2_1 _34466_ (.A(_11825_),
    .B(_11793_),
    .Y(_12115_));
 sky130_fd_sc_hd__nand2_2 _34467_ (.A(_12115_),
    .B(_11798_),
    .Y(_12116_));
 sky130_fd_sc_hd__nand3_4 _34468_ (.A(_11075_),
    .B(_11078_),
    .C(_05173_),
    .Y(_12117_));
 sky130_fd_sc_hd__o2bb2ai_4 _34469_ (.A1_N(_19575_),
    .A2_N(_07008_),
    .B1(_19923_),
    .B2(_18473_),
    .Y(_12118_));
 sky130_fd_sc_hd__o21ai_2 _34470_ (.A1(_05264_),
    .A2(_12117_),
    .B1(_12118_),
    .Y(_12119_));
 sky130_fd_sc_hd__nand2_4 _34471_ (.A(_10827_),
    .B(_05267_),
    .Y(_12120_));
 sky130_vsdinv _34472_ (.A(_12120_),
    .Y(_12121_));
 sky130_fd_sc_hd__nand2_1 _34473_ (.A(_12119_),
    .B(_12121_),
    .Y(_12122_));
 sky130_fd_sc_hd__o21ai_1 _34474_ (.A1(_19927_),
    .A2(_11762_),
    .B1(_11766_),
    .Y(_12123_));
 sky130_fd_sc_hd__nand2_2 _34475_ (.A(_12123_),
    .B(_11764_),
    .Y(_12124_));
 sky130_fd_sc_hd__o211ai_4 _34476_ (.A1(_06015_),
    .A2(_12117_),
    .B1(_12120_),
    .C1(_12118_),
    .Y(_12125_));
 sky130_fd_sc_hd__nand3_4 _34477_ (.A(_12122_),
    .B(_12124_),
    .C(_12125_),
    .Y(_12126_));
 sky130_fd_sc_hd__nand2_1 _34478_ (.A(_12119_),
    .B(_12120_),
    .Y(_12127_));
 sky130_fd_sc_hd__o211ai_4 _34479_ (.A1(_06015_),
    .A2(_12117_),
    .B1(_12121_),
    .C1(_12118_),
    .Y(_12128_));
 sky130_fd_sc_hd__nand3b_4 _34480_ (.A_N(_12124_),
    .B(_12127_),
    .C(_12128_),
    .Y(_12129_));
 sky130_fd_sc_hd__a22oi_4 _34481_ (.A1(_10835_),
    .A2(_05277_),
    .B1(\pcpi_mul.rs2[28] ),
    .B2(_19909_),
    .Y(_12130_));
 sky130_fd_sc_hd__and4_2 _34482_ (.A(_10835_),
    .B(\pcpi_mul.rs2[28] ),
    .C(_19909_),
    .D(_05277_),
    .X(_12131_));
 sky130_fd_sc_hd__nand2_2 _34483_ (.A(\pcpi_mul.rs2[27] ),
    .B(_19906_),
    .Y(_12132_));
 sky130_vsdinv _34484_ (.A(_12132_),
    .Y(_12133_));
 sky130_fd_sc_hd__o21ai_2 _34485_ (.A1(_12130_),
    .A2(_12131_),
    .B1(_12133_),
    .Y(_12134_));
 sky130_vsdinv _34486_ (.A(_12134_),
    .Y(_12135_));
 sky130_vsdinv _34487_ (.A(_12130_),
    .Y(_12136_));
 sky130_fd_sc_hd__nand3b_4 _34488_ (.A_N(_12131_),
    .B(_12136_),
    .C(_12132_),
    .Y(_12137_));
 sky130_vsdinv _34489_ (.A(_12137_),
    .Y(_12138_));
 sky130_fd_sc_hd__o2bb2ai_4 _34490_ (.A1_N(_12126_),
    .A2_N(_12129_),
    .B1(_12135_),
    .B2(_12138_),
    .Y(_12139_));
 sky130_fd_sc_hd__a21oi_2 _34491_ (.A1(_11765_),
    .A2(_11766_),
    .B1(_11774_),
    .Y(_12140_));
 sky130_fd_sc_hd__a22oi_4 _34492_ (.A1(_12140_),
    .A2(_11769_),
    .B1(_11776_),
    .B2(_11790_),
    .Y(_12141_));
 sky130_fd_sc_hd__nand2_4 _34493_ (.A(_12137_),
    .B(_12134_),
    .Y(_12142_));
 sky130_fd_sc_hd__nand3b_4 _34494_ (.A_N(_12142_),
    .B(_12129_),
    .C(_12126_),
    .Y(_12143_));
 sky130_fd_sc_hd__nand3_4 _34495_ (.A(_12139_),
    .B(_12141_),
    .C(_12143_),
    .Y(_12144_));
 sky130_fd_sc_hd__nor2_1 _34496_ (.A(_12130_),
    .B(_12131_),
    .Y(_12145_));
 sky130_fd_sc_hd__nor2_1 _34497_ (.A(_12133_),
    .B(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__or2_1 _34498_ (.A(_12130_),
    .B(_12131_),
    .X(_12147_));
 sky130_fd_sc_hd__nor2_1 _34499_ (.A(_12132_),
    .B(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__o2bb2ai_2 _34500_ (.A1_N(_12126_),
    .A2_N(_12129_),
    .B1(_12146_),
    .B2(_12148_),
    .Y(_12149_));
 sky130_fd_sc_hd__nand2_1 _34501_ (.A(_11776_),
    .B(_11790_),
    .Y(_12150_));
 sky130_fd_sc_hd__nand2_1 _34502_ (.A(_12150_),
    .B(_11771_),
    .Y(_12151_));
 sky130_fd_sc_hd__nand3_2 _34503_ (.A(_12129_),
    .B(_12126_),
    .C(_12142_),
    .Y(_12152_));
 sky130_fd_sc_hd__nand3_4 _34504_ (.A(_12149_),
    .B(_12151_),
    .C(_12152_),
    .Y(_12153_));
 sky130_fd_sc_hd__a22oi_4 _34505_ (.A1(_10256_),
    .A2(_19904_),
    .B1(_08946_),
    .B2(_06441_),
    .Y(_12154_));
 sky130_fd_sc_hd__nand3_4 _34506_ (.A(_19595_),
    .B(_08945_),
    .C(_05801_),
    .Y(_12155_));
 sky130_fd_sc_hd__nor2_4 _34507_ (.A(_06262_),
    .B(_12155_),
    .Y(_12156_));
 sky130_fd_sc_hd__nand2_4 _34508_ (.A(_19602_),
    .B(_06648_),
    .Y(_12157_));
 sky130_fd_sc_hd__o21ai_2 _34509_ (.A1(_12154_),
    .A2(_12156_),
    .B1(_12157_),
    .Y(_12158_));
 sky130_fd_sc_hd__a22o_2 _34510_ (.A1(_10256_),
    .A2(_06264_),
    .B1(_08946_),
    .B2(_07789_),
    .X(_12159_));
 sky130_vsdinv _34511_ (.A(_12157_),
    .Y(_12160_));
 sky130_fd_sc_hd__nand3b_2 _34512_ (.A_N(_12156_),
    .B(_12159_),
    .C(_12160_),
    .Y(_12161_));
 sky130_fd_sc_hd__o2111ai_4 _34513_ (.A1(_11782_),
    .A2(_11779_),
    .B1(_11786_),
    .C1(_12158_),
    .D1(_12161_),
    .Y(_12162_));
 sky130_fd_sc_hd__o21ai_4 _34514_ (.A1(_11799_),
    .A2(_11806_),
    .B1(_11808_),
    .Y(_12163_));
 sky130_fd_sc_hd__o21ai_2 _34515_ (.A1(_12154_),
    .A2(_12156_),
    .B1(_12160_),
    .Y(_12164_));
 sky130_fd_sc_hd__o21ai_2 _34516_ (.A1(_11782_),
    .A2(_11779_),
    .B1(_11786_),
    .Y(_12165_));
 sky130_fd_sc_hd__o211ai_4 _34517_ (.A1(_06829_),
    .A2(_12155_),
    .B1(_12157_),
    .C1(_12159_),
    .Y(_12166_));
 sky130_fd_sc_hd__nand3_4 _34518_ (.A(_12164_),
    .B(_12165_),
    .C(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__and3_1 _34519_ (.A(_12162_),
    .B(_12163_),
    .C(_12167_),
    .X(_12168_));
 sky130_fd_sc_hd__a21oi_4 _34520_ (.A1(_12162_),
    .A2(_12167_),
    .B1(_12163_),
    .Y(_12169_));
 sky130_fd_sc_hd__o2bb2ai_2 _34521_ (.A1_N(_12144_),
    .A2_N(_12153_),
    .B1(_12168_),
    .B2(_12169_),
    .Y(_12170_));
 sky130_fd_sc_hd__and2_1 _34522_ (.A(_12167_),
    .B(_12163_),
    .X(_12171_));
 sky130_fd_sc_hd__a21oi_4 _34523_ (.A1(_12171_),
    .A2(_12162_),
    .B1(_12169_),
    .Y(_12172_));
 sky130_fd_sc_hd__nand3_2 _34524_ (.A(_12153_),
    .B(_12172_),
    .C(_12144_),
    .Y(_12173_));
 sky130_fd_sc_hd__nand3_4 _34525_ (.A(_12116_),
    .B(_12170_),
    .C(_12173_),
    .Y(_12174_));
 sky130_fd_sc_hd__nand2_1 _34526_ (.A(_12153_),
    .B(_12144_),
    .Y(_12175_));
 sky130_fd_sc_hd__nand2_1 _34527_ (.A(_12175_),
    .B(_12172_),
    .Y(_12176_));
 sky130_fd_sc_hd__nand3b_2 _34528_ (.A_N(_12172_),
    .B(_12153_),
    .C(_12144_),
    .Y(_12177_));
 sky130_fd_sc_hd__a21oi_4 _34529_ (.A1(_11789_),
    .A2(_11791_),
    .B1(_11792_),
    .Y(_12178_));
 sky130_fd_sc_hd__a21oi_4 _34530_ (.A1(_11825_),
    .A2(_11793_),
    .B1(_12178_),
    .Y(_12179_));
 sky130_fd_sc_hd__nand3_4 _34531_ (.A(_12176_),
    .B(_12177_),
    .C(_12179_),
    .Y(_12180_));
 sky130_fd_sc_hd__a21oi_4 _34532_ (.A1(_11811_),
    .A2(_11815_),
    .B1(_11817_),
    .Y(_12181_));
 sky130_fd_sc_hd__nor2_2 _34533_ (.A(_11836_),
    .B(_11840_),
    .Y(_12182_));
 sky130_fd_sc_hd__nand2_1 _34534_ (.A(_19607_),
    .B(_06288_),
    .Y(_12183_));
 sky130_fd_sc_hd__nand3b_4 _34535_ (.A_N(_12183_),
    .B(_08541_),
    .C(_06780_),
    .Y(_12184_));
 sky130_fd_sc_hd__a22o_2 _34536_ (.A1(_08549_),
    .A2(_19894_),
    .B1(_10066_),
    .B2(_07072_),
    .X(_12185_));
 sky130_fd_sc_hd__nand2_2 _34537_ (.A(_08545_),
    .B(_19887_),
    .Y(_12186_));
 sky130_vsdinv _34538_ (.A(_12186_),
    .Y(_12187_));
 sky130_fd_sc_hd__nand3_2 _34539_ (.A(_12184_),
    .B(_12185_),
    .C(_12187_),
    .Y(_12188_));
 sky130_fd_sc_hd__a22oi_4 _34540_ (.A1(_08549_),
    .A2(_06788_),
    .B1(_08550_),
    .B2(_06462_),
    .Y(_12189_));
 sky130_fd_sc_hd__and4_2 _34541_ (.A(_10073_),
    .B(_07984_),
    .C(_06465_),
    .D(_06288_),
    .X(_12190_));
 sky130_fd_sc_hd__o21ai_2 _34542_ (.A1(_12189_),
    .A2(_12190_),
    .B1(_12186_),
    .Y(_12191_));
 sky130_fd_sc_hd__o211ai_4 _34543_ (.A1(_11834_),
    .A2(_12182_),
    .B1(_12188_),
    .C1(_12191_),
    .Y(_12192_));
 sky130_fd_sc_hd__o21ai_2 _34544_ (.A1(_12189_),
    .A2(_12190_),
    .B1(_12187_),
    .Y(_12193_));
 sky130_fd_sc_hd__a21oi_2 _34545_ (.A1(_11835_),
    .A2(_11837_),
    .B1(_11834_),
    .Y(_12194_));
 sky130_fd_sc_hd__nand3_2 _34546_ (.A(_12184_),
    .B(_12185_),
    .C(_12186_),
    .Y(_12195_));
 sky130_fd_sc_hd__nand3_4 _34547_ (.A(_12193_),
    .B(_12194_),
    .C(_12195_),
    .Y(_12196_));
 sky130_fd_sc_hd__nand2_1 _34548_ (.A(_12192_),
    .B(_12196_),
    .Y(_12197_));
 sky130_fd_sc_hd__nor2_8 _34549_ (.A(_07041_),
    .B(_07561_),
    .Y(_12198_));
 sky130_vsdinv _34550_ (.A(_12198_),
    .Y(_12199_));
 sky130_fd_sc_hd__nand2_4 _34551_ (.A(_19621_),
    .B(_06443_),
    .Y(_12200_));
 sky130_fd_sc_hd__nand2_4 _34552_ (.A(_08174_),
    .B(_06654_),
    .Y(_12201_));
 sky130_fd_sc_hd__nor2_8 _34553_ (.A(_12200_),
    .B(_12201_),
    .Y(_12202_));
 sky130_vsdinv _34554_ (.A(_12202_),
    .Y(_12203_));
 sky130_fd_sc_hd__nand2_4 _34555_ (.A(_12200_),
    .B(_12201_),
    .Y(_12204_));
 sky130_fd_sc_hd__nand3_1 _34556_ (.A(_12199_),
    .B(_12203_),
    .C(_12204_),
    .Y(_12205_));
 sky130_vsdinv _34557_ (.A(_12204_),
    .Y(_12206_));
 sky130_fd_sc_hd__o21ai_1 _34558_ (.A1(_12202_),
    .A2(_12206_),
    .B1(_12198_),
    .Y(_12207_));
 sky130_fd_sc_hd__nand2_2 _34559_ (.A(_12205_),
    .B(_12207_),
    .Y(_12208_));
 sky130_fd_sc_hd__nand2_1 _34560_ (.A(_12197_),
    .B(_12208_),
    .Y(_12209_));
 sky130_fd_sc_hd__o21ai_1 _34561_ (.A1(_12202_),
    .A2(_12206_),
    .B1(_12199_),
    .Y(_12210_));
 sky130_fd_sc_hd__nand3_1 _34562_ (.A(_12203_),
    .B(_12198_),
    .C(_12204_),
    .Y(_12211_));
 sky130_fd_sc_hd__nand2_1 _34563_ (.A(_12210_),
    .B(_12211_),
    .Y(_12212_));
 sky130_fd_sc_hd__nand3_2 _34564_ (.A(_12212_),
    .B(_12196_),
    .C(_12192_),
    .Y(_12213_));
 sky130_fd_sc_hd__nand3_4 _34565_ (.A(_12181_),
    .B(_12209_),
    .C(_12213_),
    .Y(_12214_));
 sky130_fd_sc_hd__o21ai_2 _34566_ (.A1(_11814_),
    .A2(_11823_),
    .B1(_11813_),
    .Y(_12215_));
 sky130_fd_sc_hd__nand2_1 _34567_ (.A(_12197_),
    .B(_12212_),
    .Y(_12216_));
 sky130_fd_sc_hd__nand3_4 _34568_ (.A(_12208_),
    .B(_12196_),
    .C(_12192_),
    .Y(_12217_));
 sky130_fd_sc_hd__nand3_4 _34569_ (.A(_12215_),
    .B(_12216_),
    .C(_12217_),
    .Y(_12218_));
 sky130_fd_sc_hd__nand2_1 _34570_ (.A(_12214_),
    .B(_12218_),
    .Y(_12219_));
 sky130_vsdinv _34571_ (.A(_11842_),
    .Y(_12220_));
 sky130_fd_sc_hd__a21oi_2 _34572_ (.A1(_11846_),
    .A2(_11859_),
    .B1(_12220_),
    .Y(_12221_));
 sky130_fd_sc_hd__and2_1 _34573_ (.A(_12219_),
    .B(_12221_),
    .X(_12222_));
 sky130_fd_sc_hd__a21o_1 _34574_ (.A1(_11846_),
    .A2(_11859_),
    .B1(_12220_),
    .X(_12223_));
 sky130_fd_sc_hd__and3_1 _34575_ (.A(_12214_),
    .B(_12218_),
    .C(_12223_),
    .X(_12224_));
 sky130_fd_sc_hd__o2bb2ai_4 _34576_ (.A1_N(_12174_),
    .A2_N(_12180_),
    .B1(_12222_),
    .B2(_12224_),
    .Y(_12225_));
 sky130_fd_sc_hd__clkbuf_4 _34577_ (.A(_12174_),
    .X(_12226_));
 sky130_fd_sc_hd__nand2_1 _34578_ (.A(_12219_),
    .B(_12223_),
    .Y(_12227_));
 sky130_fd_sc_hd__nand3_2 _34579_ (.A(_12214_),
    .B(_12218_),
    .C(_12221_),
    .Y(_12228_));
 sky130_fd_sc_hd__nand2_4 _34580_ (.A(_12227_),
    .B(_12228_),
    .Y(_12229_));
 sky130_fd_sc_hd__nand3_4 _34581_ (.A(_12180_),
    .B(_12226_),
    .C(_12229_),
    .Y(_12230_));
 sky130_vsdinv _34582_ (.A(_11826_),
    .Y(_12231_));
 sky130_fd_sc_hd__nand2_1 _34583_ (.A(_11820_),
    .B(_11822_),
    .Y(_12232_));
 sky130_fd_sc_hd__o2bb2ai_4 _34584_ (.A1_N(_11832_),
    .A2_N(_11878_),
    .B1(_12231_),
    .B2(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__a21oi_4 _34585_ (.A1(_12225_),
    .A2(_12230_),
    .B1(_12233_),
    .Y(_12234_));
 sky130_vsdinv _34586_ (.A(_12226_),
    .Y(_12235_));
 sky130_fd_sc_hd__nand2_2 _34587_ (.A(_12180_),
    .B(_12229_),
    .Y(_12236_));
 sky130_fd_sc_hd__o211a_1 _34588_ (.A1(_12235_),
    .A2(_12236_),
    .B1(_12225_),
    .C1(_12233_),
    .X(_12237_));
 sky130_fd_sc_hd__o22ai_4 _34589_ (.A1(_12111_),
    .A2(_12114_),
    .B1(_12234_),
    .B2(_12237_),
    .Y(_12238_));
 sky130_fd_sc_hd__o21ai_4 _34590_ (.A1(_11903_),
    .A2(_11882_),
    .B1(_11896_),
    .Y(_12239_));
 sky130_fd_sc_hd__a21oi_2 _34591_ (.A1(_12180_),
    .A2(_12226_),
    .B1(_12229_),
    .Y(_12240_));
 sky130_fd_sc_hd__and3_4 _34592_ (.A(_12180_),
    .B(_12226_),
    .C(_12229_),
    .X(_12241_));
 sky130_fd_sc_hd__a21boi_2 _34593_ (.A1(_11878_),
    .A2(_11832_),
    .B1_N(_11827_),
    .Y(_12242_));
 sky130_fd_sc_hd__o21ai_4 _34594_ (.A1(_12240_),
    .A2(_12241_),
    .B1(_12242_),
    .Y(_12243_));
 sky130_fd_sc_hd__and2_1 _34595_ (.A(_12108_),
    .B(_11718_),
    .X(_12244_));
 sky130_fd_sc_hd__a21oi_4 _34596_ (.A1(_12097_),
    .A2(_12094_),
    .B1(_12112_),
    .Y(_12245_));
 sky130_fd_sc_hd__nor2_4 _34597_ (.A(_12244_),
    .B(_12245_),
    .Y(_12246_));
 sky130_fd_sc_hd__a21oi_4 _34598_ (.A1(_12246_),
    .A2(_12113_),
    .B1(_12114_),
    .Y(_12247_));
 sky130_fd_sc_hd__nand3_4 _34599_ (.A(_12233_),
    .B(_12225_),
    .C(_12230_),
    .Y(_12248_));
 sky130_fd_sc_hd__nand3_4 _34600_ (.A(_12243_),
    .B(_12247_),
    .C(_12248_),
    .Y(_12249_));
 sky130_fd_sc_hd__nand3_4 _34601_ (.A(_12238_),
    .B(_12239_),
    .C(_12249_),
    .Y(_12250_));
 sky130_fd_sc_hd__o21ai_2 _34602_ (.A1(_12234_),
    .A2(_12237_),
    .B1(_12247_),
    .Y(_12251_));
 sky130_fd_sc_hd__a21oi_4 _34603_ (.A1(_11893_),
    .A2(_11895_),
    .B1(_11886_),
    .Y(_12252_));
 sky130_fd_sc_hd__o21ai_2 _34604_ (.A1(_12245_),
    .A2(_12098_),
    .B1(_12244_),
    .Y(_12253_));
 sky130_fd_sc_hd__o21ai_4 _34605_ (.A1(_12098_),
    .A2(_12110_),
    .B1(_12253_),
    .Y(_12254_));
 sky130_fd_sc_hd__nand3_2 _34606_ (.A(_12243_),
    .B(_12248_),
    .C(_12254_),
    .Y(_12255_));
 sky130_fd_sc_hd__nand3_4 _34607_ (.A(_12251_),
    .B(_12252_),
    .C(_12255_),
    .Y(_12256_));
 sky130_fd_sc_hd__nand2_1 _34608_ (.A(_11977_),
    .B(_11952_),
    .Y(_12257_));
 sky130_fd_sc_hd__nand2_1 _34609_ (.A(_11189_),
    .B(_11944_),
    .Y(_12258_));
 sky130_fd_sc_hd__nand2_2 _34610_ (.A(_11943_),
    .B(_12258_),
    .Y(_12259_));
 sky130_fd_sc_hd__nand2_2 _34611_ (.A(_05768_),
    .B(_10504_),
    .Y(_12260_));
 sky130_fd_sc_hd__nand2_2 _34612_ (.A(_19673_),
    .B(_19825_),
    .Y(_12261_));
 sky130_fd_sc_hd__nor2_4 _34613_ (.A(_12260_),
    .B(_12261_),
    .Y(_12262_));
 sky130_fd_sc_hd__nand2_4 _34614_ (.A(_12260_),
    .B(_12261_),
    .Y(_12263_));
 sky130_vsdinv _34615_ (.A(_12263_),
    .Y(_12264_));
 sky130_fd_sc_hd__o21ai_2 _34616_ (.A1(_12262_),
    .A2(_12264_),
    .B1(_11589_),
    .Y(_12265_));
 sky130_vsdinv _34617_ (.A(_12262_),
    .Y(_12266_));
 sky130_fd_sc_hd__nand3_2 _34618_ (.A(_12266_),
    .B(_11579_),
    .C(_12263_),
    .Y(_12267_));
 sky130_fd_sc_hd__nand3b_4 _34619_ (.A_N(_12259_),
    .B(_12265_),
    .C(_12267_),
    .Y(_12268_));
 sky130_fd_sc_hd__o21ai_2 _34620_ (.A1(_12262_),
    .A2(_12264_),
    .B1(_11579_),
    .Y(_12269_));
 sky130_fd_sc_hd__nand3_2 _34621_ (.A(_12266_),
    .B(_11589_),
    .C(_12263_),
    .Y(_12270_));
 sky130_fd_sc_hd__nand3_4 _34622_ (.A(_12269_),
    .B(_12270_),
    .C(_12259_),
    .Y(_12271_));
 sky130_fd_sc_hd__nand2_1 _34623_ (.A(_12268_),
    .B(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__o21a_2 _34624_ (.A1(_19678_),
    .A2(_19681_),
    .B1(_18467_),
    .X(_12273_));
 sky130_fd_sc_hd__buf_6 _34625_ (.A(\pcpi_mul.rs1[32] ),
    .X(_12274_));
 sky130_fd_sc_hd__nand2_4 _34626_ (.A(_12274_),
    .B(_05131_),
    .Y(_12275_));
 sky130_fd_sc_hd__a21o_1 _34627_ (.A1(_12273_),
    .A2(_11956_),
    .B1(_12275_),
    .X(_12276_));
 sky130_fd_sc_hd__nand3_4 _34628_ (.A(_12273_),
    .B(_11956_),
    .C(_12275_),
    .Y(_12277_));
 sky130_fd_sc_hd__nand2_1 _34629_ (.A(_12276_),
    .B(_12277_),
    .Y(_12278_));
 sky130_vsdinv _34630_ (.A(_12278_),
    .Y(_12279_));
 sky130_fd_sc_hd__nand2_1 _34631_ (.A(_12272_),
    .B(_12279_),
    .Y(_12280_));
 sky130_fd_sc_hd__clkbuf_2 _34632_ (.A(_12278_),
    .X(_12281_));
 sky130_fd_sc_hd__buf_2 _34633_ (.A(_12281_),
    .X(_12282_));
 sky130_fd_sc_hd__nand3_2 _34634_ (.A(_12268_),
    .B(_12271_),
    .C(_12282_),
    .Y(_12283_));
 sky130_fd_sc_hd__nand3_4 _34635_ (.A(_12257_),
    .B(_12280_),
    .C(_12283_),
    .Y(_12284_));
 sky130_fd_sc_hd__a21oi_2 _34636_ (.A1(_11963_),
    .A2(_11948_),
    .B1(_11976_),
    .Y(_12285_));
 sky130_fd_sc_hd__nand2_1 _34637_ (.A(_12272_),
    .B(_12282_),
    .Y(_12286_));
 sky130_fd_sc_hd__nand3_2 _34638_ (.A(_12268_),
    .B(_12279_),
    .C(_12271_),
    .Y(_12287_));
 sky130_fd_sc_hd__nand3_4 _34639_ (.A(_12285_),
    .B(_12286_),
    .C(_12287_),
    .Y(_12288_));
 sky130_fd_sc_hd__o21a_1 _34640_ (.A1(_11954_),
    .A2(_11955_),
    .B1(_11956_),
    .X(_12289_));
 sky130_vsdinv _34641_ (.A(_12289_),
    .Y(_12290_));
 sky130_fd_sc_hd__a21o_2 _34642_ (.A1(_12284_),
    .A2(_12288_),
    .B1(_12290_),
    .X(_12291_));
 sky130_fd_sc_hd__nand3_4 _34643_ (.A(_12284_),
    .B(_12288_),
    .C(_12290_),
    .Y(_12292_));
 sky130_fd_sc_hd__o21a_1 _34644_ (.A1(_11932_),
    .A2(_11928_),
    .B1(_11933_),
    .X(_12293_));
 sky130_fd_sc_hd__nand2_4 _34645_ (.A(_11729_),
    .B(_11740_),
    .Y(_12294_));
 sky130_fd_sc_hd__nand3_4 _34646_ (.A(_06502_),
    .B(_06488_),
    .C(_10488_),
    .Y(_12295_));
 sky130_fd_sc_hd__nor2_8 _34647_ (.A(_10497_),
    .B(_12295_),
    .Y(_12296_));
 sky130_fd_sc_hd__a22o_2 _34648_ (.A1(_19663_),
    .A2(_19844_),
    .B1(_19666_),
    .B2(_10601_),
    .X(_12297_));
 sky130_fd_sc_hd__nand2_2 _34649_ (.A(_19668_),
    .B(_10598_),
    .Y(_12298_));
 sky130_fd_sc_hd__nand3b_2 _34650_ (.A_N(_12296_),
    .B(_12297_),
    .C(_12298_),
    .Y(_12299_));
 sky130_fd_sc_hd__a21oi_2 _34651_ (.A1(_11733_),
    .A2(_11738_),
    .B1(_11737_),
    .Y(_12300_));
 sky130_fd_sc_hd__a22oi_4 _34652_ (.A1(_19663_),
    .A2(_10493_),
    .B1(_19666_),
    .B2(_11574_),
    .Y(_12301_));
 sky130_vsdinv _34653_ (.A(_12298_),
    .Y(_12302_));
 sky130_fd_sc_hd__o21ai_2 _34654_ (.A1(_12301_),
    .A2(_12296_),
    .B1(_12302_),
    .Y(_12303_));
 sky130_fd_sc_hd__nand3_4 _34655_ (.A(_12299_),
    .B(_12300_),
    .C(_12303_),
    .Y(_12304_));
 sky130_fd_sc_hd__a21o_1 _34656_ (.A1(_11733_),
    .A2(_11738_),
    .B1(_11737_),
    .X(_12305_));
 sky130_fd_sc_hd__nand3b_2 _34657_ (.A_N(_12296_),
    .B(_12297_),
    .C(_12302_),
    .Y(_12306_));
 sky130_fd_sc_hd__o21ai_2 _34658_ (.A1(_12301_),
    .A2(_12296_),
    .B1(_12298_),
    .Y(_12307_));
 sky130_fd_sc_hd__nand3_4 _34659_ (.A(_12305_),
    .B(_12306_),
    .C(_12307_),
    .Y(_12308_));
 sky130_fd_sc_hd__nor2_4 _34660_ (.A(_11912_),
    .B(_11908_),
    .Y(_12309_));
 sky130_fd_sc_hd__o2bb2ai_4 _34661_ (.A1_N(_12304_),
    .A2_N(_12308_),
    .B1(_11915_),
    .B2(_12309_),
    .Y(_12310_));
 sky130_fd_sc_hd__nor2_4 _34662_ (.A(_11915_),
    .B(_12309_),
    .Y(_12311_));
 sky130_fd_sc_hd__nand3_4 _34663_ (.A(_12308_),
    .B(_12304_),
    .C(_12311_),
    .Y(_12312_));
 sky130_fd_sc_hd__a22oi_4 _34664_ (.A1(_11728_),
    .A2(_12294_),
    .B1(_12310_),
    .B2(_12312_),
    .Y(_12313_));
 sky130_fd_sc_hd__nand2_1 _34665_ (.A(_11723_),
    .B(_11726_),
    .Y(_12314_));
 sky130_vsdinv _34666_ (.A(_12314_),
    .Y(_12315_));
 sky130_fd_sc_hd__o2111a_2 _34667_ (.A1(_11727_),
    .A2(_12315_),
    .B1(_12312_),
    .C1(_12294_),
    .D1(_12310_),
    .X(_12316_));
 sky130_vsdinv _34668_ (.A(_11917_),
    .Y(_12317_));
 sky130_fd_sc_hd__a21oi_4 _34669_ (.A1(_11922_),
    .A2(_11925_),
    .B1(_12317_),
    .Y(_12318_));
 sky130_vsdinv _34670_ (.A(_12318_),
    .Y(_12319_));
 sky130_fd_sc_hd__o21ai_2 _34671_ (.A1(_12313_),
    .A2(_12316_),
    .B1(_12319_),
    .Y(_12320_));
 sky130_fd_sc_hd__a22o_1 _34672_ (.A1(_11728_),
    .A2(_12294_),
    .B1(_12310_),
    .B2(_12312_),
    .X(_12321_));
 sky130_fd_sc_hd__o2111ai_4 _34673_ (.A1(_11727_),
    .A2(_12315_),
    .B1(_12312_),
    .C1(_12294_),
    .D1(_12310_),
    .Y(_12322_));
 sky130_fd_sc_hd__nand3_2 _34674_ (.A(_12321_),
    .B(_12322_),
    .C(_12318_),
    .Y(_12323_));
 sky130_fd_sc_hd__nand3_4 _34675_ (.A(_12293_),
    .B(_12320_),
    .C(_12323_),
    .Y(_12324_));
 sky130_fd_sc_hd__o21ai_2 _34676_ (.A1(_12313_),
    .A2(_12316_),
    .B1(_12318_),
    .Y(_12325_));
 sky130_fd_sc_hd__o21ai_2 _34677_ (.A1(_11932_),
    .A2(_11928_),
    .B1(_11933_),
    .Y(_12326_));
 sky130_fd_sc_hd__nand3_2 _34678_ (.A(_12321_),
    .B(_12319_),
    .C(_12322_),
    .Y(_12327_));
 sky130_fd_sc_hd__nand3_4 _34679_ (.A(_12325_),
    .B(_12326_),
    .C(_12327_),
    .Y(_12328_));
 sky130_fd_sc_hd__a22oi_4 _34680_ (.A1(_12291_),
    .A2(_12292_),
    .B1(_12324_),
    .B2(_12328_),
    .Y(_12329_));
 sky130_vsdinv _34681_ (.A(_12288_),
    .Y(_12330_));
 sky130_fd_sc_hd__nand2_2 _34682_ (.A(_12284_),
    .B(_12290_),
    .Y(_12331_));
 sky130_fd_sc_hd__o2111a_1 _34683_ (.A1(_12330_),
    .A2(_12331_),
    .B1(_12291_),
    .C1(_12328_),
    .D1(_12324_),
    .X(_12332_));
 sky130_vsdinv _34684_ (.A(_11747_),
    .Y(_12333_));
 sky130_fd_sc_hd__nand2_1 _34685_ (.A(_11745_),
    .B(_11746_),
    .Y(_12334_));
 sky130_fd_sc_hd__o2bb2ai_4 _34686_ (.A1_N(_11757_),
    .A2_N(_11760_),
    .B1(_12333_),
    .B2(_12334_),
    .Y(_12335_));
 sky130_fd_sc_hd__o21bai_4 _34687_ (.A1(_12329_),
    .A2(_12332_),
    .B1_N(_12335_),
    .Y(_12336_));
 sky130_fd_sc_hd__a22o_1 _34688_ (.A1(_12291_),
    .A2(_12292_),
    .B1(_12324_),
    .B2(_12328_),
    .X(_12337_));
 sky130_fd_sc_hd__o2111ai_4 _34689_ (.A1(_12330_),
    .A2(_12331_),
    .B1(_12291_),
    .C1(_12328_),
    .D1(_12324_),
    .Y(_12338_));
 sky130_fd_sc_hd__nand3_4 _34690_ (.A(_12337_),
    .B(_12338_),
    .C(_12335_),
    .Y(_12339_));
 sky130_vsdinv _34691_ (.A(_11940_),
    .Y(_12340_));
 sky130_fd_sc_hd__a21oi_4 _34692_ (.A1(_11936_),
    .A2(_11981_),
    .B1(_12340_),
    .Y(_12341_));
 sky130_vsdinv _34693_ (.A(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__a21oi_4 _34694_ (.A1(_12336_),
    .A2(_12339_),
    .B1(_12342_),
    .Y(_12343_));
 sky130_fd_sc_hd__nand3_2 _34695_ (.A(_12342_),
    .B(_12336_),
    .C(_12339_),
    .Y(_12344_));
 sky130_vsdinv _34696_ (.A(_12344_),
    .Y(_12345_));
 sky130_fd_sc_hd__o2bb2ai_4 _34697_ (.A1_N(_12250_),
    .A2_N(_12256_),
    .B1(_12343_),
    .B2(_12345_),
    .Y(_12346_));
 sky130_fd_sc_hd__nand2_1 _34698_ (.A(_12337_),
    .B(_12338_),
    .Y(_12347_));
 sky130_vsdinv _34699_ (.A(_12335_),
    .Y(_12348_));
 sky130_fd_sc_hd__a21oi_4 _34700_ (.A1(_12347_),
    .A2(_12348_),
    .B1(_12341_),
    .Y(_12349_));
 sky130_fd_sc_hd__a21oi_4 _34701_ (.A1(_12339_),
    .A2(_12349_),
    .B1(_12343_),
    .Y(_12350_));
 sky130_fd_sc_hd__nand3_4 _34702_ (.A(_12350_),
    .B(_12250_),
    .C(_12256_),
    .Y(_12351_));
 sky130_fd_sc_hd__nand2_1 _34703_ (.A(_12005_),
    .B(_11905_),
    .Y(_12352_));
 sky130_fd_sc_hd__nand2_4 _34704_ (.A(_12352_),
    .B(_11898_),
    .Y(_12353_));
 sky130_fd_sc_hd__a21oi_4 _34705_ (.A1(_12346_),
    .A2(_12351_),
    .B1(_12353_),
    .Y(_12354_));
 sky130_vsdinv _34706_ (.A(_11898_),
    .Y(_12355_));
 sky130_fd_sc_hd__a32oi_2 _34707_ (.A1(_11899_),
    .A2(_11900_),
    .A3(_11904_),
    .B1(_12002_),
    .B2(_12004_),
    .Y(_12356_));
 sky130_fd_sc_hd__o211a_2 _34708_ (.A1(_12355_),
    .A2(_12356_),
    .B1(_12351_),
    .C1(_12346_),
    .X(_12357_));
 sky130_fd_sc_hd__nor2_4 _34709_ (.A(_11978_),
    .B(_11987_),
    .Y(_12358_));
 sky130_fd_sc_hd__and3_2 _34710_ (.A(_11997_),
    .B(_11992_),
    .C(_12358_),
    .X(_12359_));
 sky130_fd_sc_hd__and2_1 _34711_ (.A(_11997_),
    .B(_11992_),
    .X(_12360_));
 sky130_fd_sc_hd__nor2_2 _34712_ (.A(_12358_),
    .B(_12360_),
    .Y(_12361_));
 sky130_fd_sc_hd__nor2_4 _34713_ (.A(_12359_),
    .B(_12361_),
    .Y(_12362_));
 sky130_fd_sc_hd__o21ai_2 _34714_ (.A1(_12354_),
    .A2(_12357_),
    .B1(_12362_),
    .Y(_12363_));
 sky130_fd_sc_hd__a21oi_4 _34715_ (.A1(_12017_),
    .A2(_12026_),
    .B1(_12011_),
    .Y(_12364_));
 sky130_fd_sc_hd__a21o_1 _34716_ (.A1(_12346_),
    .A2(_12351_),
    .B1(_12353_),
    .X(_12365_));
 sky130_fd_sc_hd__nand3_4 _34717_ (.A(_12353_),
    .B(_12351_),
    .C(_12346_),
    .Y(_12366_));
 sky130_fd_sc_hd__xnor2_2 _34718_ (.A(_12358_),
    .B(_12360_),
    .Y(_12367_));
 sky130_fd_sc_hd__nand3_2 _34719_ (.A(_12365_),
    .B(_12366_),
    .C(_12367_),
    .Y(_12368_));
 sky130_fd_sc_hd__nand3_4 _34720_ (.A(_12363_),
    .B(_12364_),
    .C(_12368_),
    .Y(_12369_));
 sky130_fd_sc_hd__buf_2 _34721_ (.A(_12361_),
    .X(_12370_));
 sky130_fd_sc_hd__o22ai_4 _34722_ (.A1(_12370_),
    .A2(_12359_),
    .B1(_12354_),
    .B2(_12357_),
    .Y(_12371_));
 sky130_fd_sc_hd__nand3_2 _34723_ (.A(_12365_),
    .B(_12366_),
    .C(_12362_),
    .Y(_12372_));
 sky130_fd_sc_hd__o21ai_2 _34724_ (.A1(_12019_),
    .A2(_12009_),
    .B1(_12018_),
    .Y(_12373_));
 sky130_fd_sc_hd__nand3_4 _34725_ (.A(_12371_),
    .B(_12372_),
    .C(_12373_),
    .Y(_12374_));
 sky130_fd_sc_hd__nand3_2 _34726_ (.A(_12369_),
    .B(_12374_),
    .C(_12022_),
    .Y(_12375_));
 sky130_vsdinv _34727_ (.A(_12375_),
    .Y(_12376_));
 sky130_vsdinv _34728_ (.A(_12022_),
    .Y(_12377_));
 sky130_fd_sc_hd__nand2_1 _34729_ (.A(_12369_),
    .B(_12374_),
    .Y(_12378_));
 sky130_fd_sc_hd__a31oi_2 _34730_ (.A1(_11683_),
    .A2(_12012_),
    .A3(_12020_),
    .B1(_11658_),
    .Y(_12379_));
 sky130_fd_sc_hd__o2bb2ai_2 _34731_ (.A1_N(_12377_),
    .A2_N(_12378_),
    .B1(_12035_),
    .B2(_12379_),
    .Y(_12380_));
 sky130_fd_sc_hd__o2bb2ai_1 _34732_ (.A1_N(_12374_),
    .A2_N(_12369_),
    .B1(_11689_),
    .B2(_11687_),
    .Y(_12381_));
 sky130_fd_sc_hd__nand2_1 _34733_ (.A(_12036_),
    .B(_12028_),
    .Y(_12382_));
 sky130_fd_sc_hd__a21o_1 _34734_ (.A1(_12381_),
    .A2(_12375_),
    .B1(_12382_),
    .X(_12383_));
 sky130_fd_sc_hd__o21a_2 _34735_ (.A1(_12376_),
    .A2(_12380_),
    .B1(_12383_),
    .X(_12384_));
 sky130_fd_sc_hd__nand2_1 _34736_ (.A(_12042_),
    .B(_12038_),
    .Y(_12385_));
 sky130_fd_sc_hd__nand2_2 _34737_ (.A(_12385_),
    .B(_12034_),
    .Y(_12386_));
 sky130_fd_sc_hd__xnor2_4 _34738_ (.A(_12384_),
    .B(_12386_),
    .Y(_02654_));
 sky130_fd_sc_hd__a21oi_4 _34739_ (.A1(_12365_),
    .A2(_12362_),
    .B1(_12357_),
    .Y(_12387_));
 sky130_fd_sc_hd__nand2_2 _34740_ (.A(_12233_),
    .B(_12225_),
    .Y(_12388_));
 sky130_fd_sc_hd__o22ai_4 _34741_ (.A1(_12241_),
    .A2(_12388_),
    .B1(_12254_),
    .B2(_12234_),
    .Y(_12389_));
 sky130_fd_sc_hd__nand2_1 _34742_ (.A(_12236_),
    .B(_12226_),
    .Y(_12390_));
 sky130_fd_sc_hd__nand2_2 _34743_ (.A(_12172_),
    .B(_12144_),
    .Y(_12391_));
 sky130_fd_sc_hd__nand2_2 _34744_ (.A(_12391_),
    .B(_12153_),
    .Y(_12392_));
 sky130_fd_sc_hd__nand3_4 _34745_ (.A(_11080_),
    .B(_19575_),
    .C(_05208_),
    .Y(_12393_));
 sky130_fd_sc_hd__nand2_1 _34746_ (.A(_19575_),
    .B(_05377_),
    .Y(_12394_));
 sky130_fd_sc_hd__o21ai_4 _34747_ (.A1(_05224_),
    .A2(_18473_),
    .B1(_12394_),
    .Y(_12395_));
 sky130_fd_sc_hd__o21ai_2 _34748_ (.A1(_06330_),
    .A2(_12393_),
    .B1(_12395_),
    .Y(_12396_));
 sky130_fd_sc_hd__nand2_4 _34749_ (.A(_10827_),
    .B(_05379_),
    .Y(_12397_));
 sky130_fd_sc_hd__nand2_1 _34750_ (.A(_12396_),
    .B(_12397_),
    .Y(_12398_));
 sky130_vsdinv _34751_ (.A(_12397_),
    .Y(_12399_));
 sky130_fd_sc_hd__o211ai_4 _34752_ (.A1(_05237_),
    .A2(_12393_),
    .B1(_12399_),
    .C1(_12395_),
    .Y(_12400_));
 sky130_fd_sc_hd__buf_6 _34753_ (.A(_19575_),
    .X(_12401_));
 sky130_fd_sc_hd__buf_8 _34754_ (.A(_11080_),
    .X(_12402_));
 sky130_fd_sc_hd__a22oi_4 _34755_ (.A1(_12401_),
    .A2(_06330_),
    .B1(_05154_),
    .B2(_12402_),
    .Y(_12403_));
 sky130_fd_sc_hd__o22ai_4 _34756_ (.A1(_06015_),
    .A2(_12117_),
    .B1(_12120_),
    .B2(_12403_),
    .Y(_12404_));
 sky130_fd_sc_hd__nand3_4 _34757_ (.A(_12398_),
    .B(_12400_),
    .C(_12404_),
    .Y(_12405_));
 sky130_fd_sc_hd__nand2_1 _34758_ (.A(_12396_),
    .B(_12399_),
    .Y(_12406_));
 sky130_fd_sc_hd__o21ai_1 _34759_ (.A1(_05147_),
    .A2(_12117_),
    .B1(_12120_),
    .Y(_12407_));
 sky130_fd_sc_hd__nand2_2 _34760_ (.A(_12407_),
    .B(_12118_),
    .Y(_12408_));
 sky130_fd_sc_hd__o211ai_4 _34761_ (.A1(_19921_),
    .A2(_12393_),
    .B1(_12397_),
    .C1(_12395_),
    .Y(_12409_));
 sky130_fd_sc_hd__nand3_4 _34762_ (.A(_12406_),
    .B(_12408_),
    .C(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__a22oi_4 _34763_ (.A1(_10836_),
    .A2(_19910_),
    .B1(net494),
    .B2(_05661_),
    .Y(_12411_));
 sky130_fd_sc_hd__nand2_2 _34764_ (.A(_19582_),
    .B(_05488_),
    .Y(_12412_));
 sky130_fd_sc_hd__nand2_2 _34765_ (.A(_10046_),
    .B(_06105_),
    .Y(_12413_));
 sky130_fd_sc_hd__nor2_4 _34766_ (.A(_12412_),
    .B(_12413_),
    .Y(_12414_));
 sky130_fd_sc_hd__nand2_2 _34767_ (.A(_19591_),
    .B(_05796_),
    .Y(_12415_));
 sky130_vsdinv _34768_ (.A(_12415_),
    .Y(_12416_));
 sky130_fd_sc_hd__o21ai_1 _34769_ (.A1(_12411_),
    .A2(_12414_),
    .B1(_12416_),
    .Y(_12417_));
 sky130_vsdinv _34770_ (.A(_12417_),
    .Y(_12418_));
 sky130_fd_sc_hd__nand3b_4 _34771_ (.A_N(_12412_),
    .B(_10282_),
    .C(_06686_),
    .Y(_12419_));
 sky130_fd_sc_hd__nand2_2 _34772_ (.A(_12412_),
    .B(_12413_),
    .Y(_12420_));
 sky130_fd_sc_hd__nand3_2 _34773_ (.A(_12419_),
    .B(_12415_),
    .C(_12420_),
    .Y(_12421_));
 sky130_vsdinv _34774_ (.A(_12421_),
    .Y(_12422_));
 sky130_fd_sc_hd__o2bb2ai_2 _34775_ (.A1_N(_12405_),
    .A2_N(_12410_),
    .B1(_12418_),
    .B2(_12422_),
    .Y(_12423_));
 sky130_fd_sc_hd__a21oi_2 _34776_ (.A1(_12119_),
    .A2(_12120_),
    .B1(_12124_),
    .Y(_12424_));
 sky130_fd_sc_hd__a22oi_4 _34777_ (.A1(_12424_),
    .A2(_12128_),
    .B1(_12126_),
    .B2(_12142_),
    .Y(_12425_));
 sky130_fd_sc_hd__nand2_2 _34778_ (.A(_12417_),
    .B(_12421_),
    .Y(_12426_));
 sky130_fd_sc_hd__nand3b_2 _34779_ (.A_N(_12426_),
    .B(_12405_),
    .C(_12410_),
    .Y(_12427_));
 sky130_fd_sc_hd__nand3_4 _34780_ (.A(_12423_),
    .B(_12425_),
    .C(_12427_),
    .Y(_12428_));
 sky130_fd_sc_hd__nand2_1 _34781_ (.A(_12126_),
    .B(_12142_),
    .Y(_12429_));
 sky130_fd_sc_hd__nand2_2 _34782_ (.A(_12429_),
    .B(_12129_),
    .Y(_12430_));
 sky130_fd_sc_hd__nor2_1 _34783_ (.A(_12411_),
    .B(_12414_),
    .Y(_12431_));
 sky130_fd_sc_hd__nor2_1 _34784_ (.A(_12416_),
    .B(_12431_),
    .Y(_12432_));
 sky130_fd_sc_hd__and3_1 _34785_ (.A(_12419_),
    .B(_12416_),
    .C(_12420_),
    .X(_12433_));
 sky130_fd_sc_hd__o2bb2ai_1 _34786_ (.A1_N(_12405_),
    .A2_N(_12410_),
    .B1(_12432_),
    .B2(_12433_),
    .Y(_12434_));
 sky130_fd_sc_hd__nand3_2 _34787_ (.A(_12405_),
    .B(_12410_),
    .C(_12426_),
    .Y(_12435_));
 sky130_fd_sc_hd__nand3_4 _34788_ (.A(_12430_),
    .B(_12434_),
    .C(_12435_),
    .Y(_12436_));
 sky130_fd_sc_hd__o21a_1 _34789_ (.A1(_12133_),
    .A2(_12131_),
    .B1(_12136_),
    .X(_12437_));
 sky130_fd_sc_hd__nand3_4 _34790_ (.A(_19596_),
    .B(_09227_),
    .C(_06448_),
    .Y(_12438_));
 sky130_fd_sc_hd__nor2_4 _34791_ (.A(_05787_),
    .B(_12438_),
    .Y(_12439_));
 sky130_fd_sc_hd__a22o_2 _34792_ (.A1(_10260_),
    .A2(_05804_),
    .B1(_09723_),
    .B2(_05977_),
    .X(_12440_));
 sky130_fd_sc_hd__nand2_2 _34793_ (.A(_11801_),
    .B(_06652_),
    .Y(_12441_));
 sky130_vsdinv _34794_ (.A(_12441_),
    .Y(_12442_));
 sky130_fd_sc_hd__nand3b_4 _34795_ (.A_N(_12439_),
    .B(_12440_),
    .C(_12442_),
    .Y(_12443_));
 sky130_fd_sc_hd__a22oi_4 _34796_ (.A1(_09485_),
    .A2(_06260_),
    .B1(_10261_),
    .B2(_05977_),
    .Y(_12444_));
 sky130_fd_sc_hd__o21ai_2 _34797_ (.A1(_12444_),
    .A2(_12439_),
    .B1(_12441_),
    .Y(_12445_));
 sky130_fd_sc_hd__nand3_4 _34798_ (.A(_12437_),
    .B(_12443_),
    .C(_12445_),
    .Y(_12446_));
 sky130_fd_sc_hd__o21ai_2 _34799_ (.A1(_12133_),
    .A2(_12131_),
    .B1(_12136_),
    .Y(_12447_));
 sky130_fd_sc_hd__o21ai_2 _34800_ (.A1(_12444_),
    .A2(_12439_),
    .B1(_12442_),
    .Y(_12448_));
 sky130_fd_sc_hd__o211ai_4 _34801_ (.A1(_07102_),
    .A2(_12438_),
    .B1(_12441_),
    .C1(_12440_),
    .Y(_12449_));
 sky130_fd_sc_hd__nand3_4 _34802_ (.A(_12447_),
    .B(_12448_),
    .C(_12449_),
    .Y(_12450_));
 sky130_fd_sc_hd__a21o_2 _34803_ (.A1(_12159_),
    .A2(_12160_),
    .B1(_12156_),
    .X(_12451_));
 sky130_fd_sc_hd__and3_1 _34804_ (.A(_12446_),
    .B(_12450_),
    .C(_12451_),
    .X(_12452_));
 sky130_fd_sc_hd__a21oi_4 _34805_ (.A1(_12446_),
    .A2(_12450_),
    .B1(_12451_),
    .Y(_12453_));
 sky130_fd_sc_hd__o2bb2ai_4 _34806_ (.A1_N(_12428_),
    .A2_N(_12436_),
    .B1(_12452_),
    .B2(_12453_),
    .Y(_12454_));
 sky130_fd_sc_hd__and2_1 _34807_ (.A(_12450_),
    .B(_12451_),
    .X(_12455_));
 sky130_fd_sc_hd__a21oi_4 _34808_ (.A1(_12455_),
    .A2(_12446_),
    .B1(_12453_),
    .Y(_12456_));
 sky130_fd_sc_hd__nand3_4 _34809_ (.A(_12456_),
    .B(_12436_),
    .C(_12428_),
    .Y(_12457_));
 sky130_fd_sc_hd__nand3_4 _34810_ (.A(_12392_),
    .B(_12454_),
    .C(_12457_),
    .Y(_12458_));
 sky130_fd_sc_hd__nand2_2 _34811_ (.A(_12436_),
    .B(_12428_),
    .Y(_12459_));
 sky130_fd_sc_hd__nand2_1 _34812_ (.A(_12459_),
    .B(_12456_),
    .Y(_12460_));
 sky130_fd_sc_hd__a21oi_4 _34813_ (.A1(_12139_),
    .A2(_12143_),
    .B1(_12141_),
    .Y(_12461_));
 sky130_fd_sc_hd__a21oi_2 _34814_ (.A1(_12144_),
    .A2(_12172_),
    .B1(_12461_),
    .Y(_12462_));
 sky130_fd_sc_hd__a21o_1 _34815_ (.A1(_12455_),
    .A2(_12446_),
    .B1(_12453_),
    .X(_12463_));
 sky130_fd_sc_hd__nand3_2 _34816_ (.A(_12463_),
    .B(_12428_),
    .C(_12436_),
    .Y(_12464_));
 sky130_fd_sc_hd__nand3_4 _34817_ (.A(_12460_),
    .B(_12462_),
    .C(_12464_),
    .Y(_12465_));
 sky130_fd_sc_hd__buf_6 _34818_ (.A(_10066_),
    .X(_12466_));
 sky130_fd_sc_hd__a22oi_4 _34819_ (.A1(_19608_),
    .A2(_06284_),
    .B1(_12466_),
    .B2(_11848_),
    .Y(_12467_));
 sky130_fd_sc_hd__buf_4 _34820_ (.A(_08152_),
    .X(_12468_));
 sky130_fd_sc_hd__and4_2 _34821_ (.A(_12468_),
    .B(_08155_),
    .C(_07327_),
    .D(_06286_),
    .X(_12469_));
 sky130_fd_sc_hd__buf_4 _34822_ (.A(_08545_),
    .X(_12470_));
 sky130_fd_sc_hd__nand2_2 _34823_ (.A(_12470_),
    .B(_19884_),
    .Y(_12471_));
 sky130_vsdinv _34824_ (.A(_12471_),
    .Y(_12472_));
 sky130_fd_sc_hd__o21ai_2 _34825_ (.A1(_12467_),
    .A2(_12469_),
    .B1(_12472_),
    .Y(_12473_));
 sky130_fd_sc_hd__a21oi_4 _34826_ (.A1(_12185_),
    .A2(_12187_),
    .B1(_12190_),
    .Y(_12474_));
 sky130_fd_sc_hd__nand2_1 _34827_ (.A(_12468_),
    .B(_06780_),
    .Y(_12475_));
 sky130_fd_sc_hd__nand3b_4 _34828_ (.A_N(_12475_),
    .B(_12466_),
    .C(net435),
    .Y(_12476_));
 sky130_fd_sc_hd__a22o_1 _34829_ (.A1(_12468_),
    .A2(_06284_),
    .B1(_19612_),
    .B2(_06640_),
    .X(_12477_));
 sky130_fd_sc_hd__nand3_2 _34830_ (.A(_12476_),
    .B(_12471_),
    .C(_12477_),
    .Y(_12478_));
 sky130_fd_sc_hd__nand3_4 _34831_ (.A(_12473_),
    .B(_12474_),
    .C(_12478_),
    .Y(_12479_));
 sky130_vsdinv _34832_ (.A(_12479_),
    .Y(_12480_));
 sky130_fd_sc_hd__a22oi_4 _34833_ (.A1(_11847_),
    .A2(_07055_),
    .B1(_11849_),
    .B2(_07344_),
    .Y(_12481_));
 sky130_fd_sc_hd__nand2_2 _34834_ (.A(_07934_),
    .B(_07052_),
    .Y(_12482_));
 sky130_fd_sc_hd__nand2_2 _34835_ (.A(_07825_),
    .B(_08734_),
    .Y(_12483_));
 sky130_fd_sc_hd__nor2_4 _34836_ (.A(_12482_),
    .B(_12483_),
    .Y(_12484_));
 sky130_fd_sc_hd__nor2_1 _34837_ (.A(_12481_),
    .B(_12484_),
    .Y(_12485_));
 sky130_fd_sc_hd__nor2_4 _34838_ (.A(net471),
    .B(_10724_),
    .Y(_12486_));
 sky130_vsdinv _34839_ (.A(_12486_),
    .Y(_12487_));
 sky130_fd_sc_hd__nand2_1 _34840_ (.A(_12485_),
    .B(_12487_),
    .Y(_12488_));
 sky130_fd_sc_hd__o21ai_2 _34841_ (.A1(_12481_),
    .A2(_12484_),
    .B1(_12486_),
    .Y(_12489_));
 sky130_fd_sc_hd__nand2_4 _34842_ (.A(_12488_),
    .B(_12489_),
    .Y(_12490_));
 sky130_fd_sc_hd__o21ai_2 _34843_ (.A1(_12467_),
    .A2(_12469_),
    .B1(_12471_),
    .Y(_12491_));
 sky130_fd_sc_hd__nand3_2 _34844_ (.A(_12476_),
    .B(_12472_),
    .C(_12477_),
    .Y(_12492_));
 sky130_fd_sc_hd__o21ai_2 _34845_ (.A1(_12186_),
    .A2(_12189_),
    .B1(_12184_),
    .Y(_12493_));
 sky130_fd_sc_hd__nand3_4 _34846_ (.A(_12491_),
    .B(_12492_),
    .C(_12493_),
    .Y(_12494_));
 sky130_fd_sc_hd__nand2_1 _34847_ (.A(_12490_),
    .B(_12494_),
    .Y(_12495_));
 sky130_fd_sc_hd__nand2_1 _34848_ (.A(_12167_),
    .B(_12163_),
    .Y(_12496_));
 sky130_fd_sc_hd__nand2_2 _34849_ (.A(_12496_),
    .B(_12162_),
    .Y(_12497_));
 sky130_fd_sc_hd__a21o_2 _34850_ (.A1(_12479_),
    .A2(_12494_),
    .B1(_12490_),
    .X(_12498_));
 sky130_fd_sc_hd__o211a_2 _34851_ (.A1(_12480_),
    .A2(_12495_),
    .B1(_12497_),
    .C1(_12498_),
    .X(_12499_));
 sky130_fd_sc_hd__nand3_4 _34852_ (.A(_12490_),
    .B(_12479_),
    .C(_12494_),
    .Y(_12500_));
 sky130_vsdinv _34853_ (.A(_12167_),
    .Y(_12501_));
 sky130_fd_sc_hd__and2b_1 _34854_ (.A_N(_12163_),
    .B(_12162_),
    .X(_12502_));
 sky130_fd_sc_hd__o2bb2ai_4 _34855_ (.A1_N(_12500_),
    .A2_N(_12498_),
    .B1(_12501_),
    .B2(_12502_),
    .Y(_12503_));
 sky130_fd_sc_hd__nand2_4 _34856_ (.A(_12217_),
    .B(_12192_),
    .Y(_12504_));
 sky130_fd_sc_hd__nand2_2 _34857_ (.A(_12503_),
    .B(_12504_),
    .Y(_12505_));
 sky130_fd_sc_hd__nor2_1 _34858_ (.A(_12499_),
    .B(_12505_),
    .Y(_12506_));
 sky130_fd_sc_hd__nand3_4 _34859_ (.A(_12498_),
    .B(_12497_),
    .C(_12500_),
    .Y(_12507_));
 sky130_fd_sc_hd__a21oi_4 _34860_ (.A1(_12503_),
    .A2(_12507_),
    .B1(_12504_),
    .Y(_12508_));
 sky130_fd_sc_hd__o2bb2ai_2 _34861_ (.A1_N(_12458_),
    .A2_N(_12465_),
    .B1(_12506_),
    .B2(_12508_),
    .Y(_12509_));
 sky130_fd_sc_hd__and2_2 _34862_ (.A(_12217_),
    .B(_12192_),
    .X(_12510_));
 sky130_fd_sc_hd__a21oi_4 _34863_ (.A1(_12498_),
    .A2(_12500_),
    .B1(_12497_),
    .Y(_12511_));
 sky130_fd_sc_hd__nor2_2 _34864_ (.A(_12510_),
    .B(_12511_),
    .Y(_12512_));
 sky130_fd_sc_hd__a21oi_4 _34865_ (.A1(_12507_),
    .A2(_12512_),
    .B1(_12508_),
    .Y(_12513_));
 sky130_fd_sc_hd__nand3_4 _34866_ (.A(_12513_),
    .B(_12465_),
    .C(_12458_),
    .Y(_12514_));
 sky130_fd_sc_hd__nand3_4 _34867_ (.A(_12390_),
    .B(_12509_),
    .C(_12514_),
    .Y(_12515_));
 sky130_fd_sc_hd__nand2_2 _34868_ (.A(_12465_),
    .B(_12458_),
    .Y(_12516_));
 sky130_fd_sc_hd__nand2_1 _34869_ (.A(_12516_),
    .B(_12513_),
    .Y(_12517_));
 sky130_fd_sc_hd__a21boi_4 _34870_ (.A1(_12180_),
    .A2(_12229_),
    .B1_N(_12174_),
    .Y(_12518_));
 sky130_fd_sc_hd__o21ai_2 _34871_ (.A1(_12511_),
    .A2(_12499_),
    .B1(_12510_),
    .Y(_12519_));
 sky130_fd_sc_hd__o21ai_4 _34872_ (.A1(_12499_),
    .A2(_12505_),
    .B1(_12519_),
    .Y(_12520_));
 sky130_fd_sc_hd__nand3_2 _34873_ (.A(_12520_),
    .B(_12465_),
    .C(_12458_),
    .Y(_12521_));
 sky130_fd_sc_hd__nand3_4 _34874_ (.A(_12517_),
    .B(_12518_),
    .C(_12521_),
    .Y(_12522_));
 sky130_fd_sc_hd__nand3_4 _34875_ (.A(_07007_),
    .B(_06897_),
    .C(_19861_),
    .Y(_12523_));
 sky130_fd_sc_hd__a22o_4 _34876_ (.A1(_07007_),
    .A2(_19861_),
    .B1(_06906_),
    .B2(_09972_),
    .X(_12524_));
 sky130_fd_sc_hd__o21ai_2 _34877_ (.A1(_10466_),
    .A2(_12523_),
    .B1(_12524_),
    .Y(_12525_));
 sky130_fd_sc_hd__o21ai_4 _34878_ (.A1(_11721_),
    .A2(_10652_),
    .B1(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__nor2_4 _34879_ (.A(_10449_),
    .B(_12523_),
    .Y(_12527_));
 sky130_fd_sc_hd__nor2_8 _34880_ (.A(_06030_),
    .B(_09806_),
    .Y(_12528_));
 sky130_fd_sc_hd__nand3b_4 _34881_ (.A_N(_12527_),
    .B(_12524_),
    .C(_12528_),
    .Y(_12529_));
 sky130_fd_sc_hd__a21o_2 _34882_ (.A1(_12069_),
    .A2(_12071_),
    .B1(_12068_),
    .X(_12530_));
 sky130_fd_sc_hd__a21o_2 _34883_ (.A1(_12526_),
    .A2(_12529_),
    .B1(_12530_),
    .X(_12531_));
 sky130_fd_sc_hd__nand3_4 _34884_ (.A(_12526_),
    .B(_12530_),
    .C(_12529_),
    .Y(_12532_));
 sky130_fd_sc_hd__a22oi_4 _34885_ (.A1(_06156_),
    .A2(_09075_),
    .B1(_05883_),
    .B2(_11228_),
    .Y(_12533_));
 sky130_fd_sc_hd__and4_1 _34886_ (.A(_06401_),
    .B(_06158_),
    .C(_19847_),
    .D(_09079_),
    .X(_12534_));
 sky130_fd_sc_hd__buf_2 _34887_ (.A(_12534_),
    .X(_12535_));
 sky130_fd_sc_hd__nor2_1 _34888_ (.A(_12533_),
    .B(_12535_),
    .Y(_12536_));
 sky130_fd_sc_hd__nand2_2 _34889_ (.A(_05731_),
    .B(_09947_),
    .Y(_12537_));
 sky130_fd_sc_hd__nand2_1 _34890_ (.A(_12536_),
    .B(_12537_),
    .Y(_12538_));
 sky130_vsdinv _34891_ (.A(_12537_),
    .Y(_12539_));
 sky130_fd_sc_hd__o21ai_2 _34892_ (.A1(_12533_),
    .A2(_12535_),
    .B1(_12539_),
    .Y(_12540_));
 sky130_fd_sc_hd__nand2_4 _34893_ (.A(_12538_),
    .B(_12540_),
    .Y(_12541_));
 sky130_fd_sc_hd__a21oi_4 _34894_ (.A1(_12531_),
    .A2(_12532_),
    .B1(_12541_),
    .Y(_12542_));
 sky130_fd_sc_hd__and3_1 _34895_ (.A(_12526_),
    .B(_12530_),
    .C(_12529_),
    .X(_12543_));
 sky130_fd_sc_hd__buf_2 _34896_ (.A(_12543_),
    .X(_12544_));
 sky130_fd_sc_hd__nand2_2 _34897_ (.A(_12531_),
    .B(_12541_),
    .Y(_12545_));
 sky130_fd_sc_hd__nor2_2 _34898_ (.A(_12544_),
    .B(_12545_),
    .Y(_12546_));
 sky130_fd_sc_hd__a31o_1 _34899_ (.A1(_12204_),
    .A2(_11003_),
    .A3(_19879_),
    .B1(_12202_),
    .X(_12547_));
 sky130_fd_sc_hd__nand2_1 _34900_ (.A(_11695_),
    .B(_10394_),
    .Y(_12548_));
 sky130_fd_sc_hd__nand3b_4 _34901_ (.A_N(_12548_),
    .B(_10999_),
    .C(_19869_),
    .Y(_12549_));
 sky130_fd_sc_hd__nand2_4 _34902_ (.A(_19641_),
    .B(_08333_),
    .Y(_12550_));
 sky130_vsdinv _34903_ (.A(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__a22o_2 _34904_ (.A1(_19632_),
    .A2(_19871_),
    .B1(_19636_),
    .B2(_10149_),
    .X(_12552_));
 sky130_fd_sc_hd__nand3_4 _34905_ (.A(_12549_),
    .B(_12551_),
    .C(_12552_),
    .Y(_12553_));
 sky130_fd_sc_hd__a22oi_4 _34906_ (.A1(_11695_),
    .A2(_10394_),
    .B1(_08873_),
    .B2(_10395_),
    .Y(_12554_));
 sky130_fd_sc_hd__and4_2 _34907_ (.A(_11695_),
    .B(_08623_),
    .C(_10395_),
    .D(_10394_),
    .X(_12555_));
 sky130_fd_sc_hd__o21ai_2 _34908_ (.A1(_12554_),
    .A2(_12555_),
    .B1(_12550_),
    .Y(_12556_));
 sky130_fd_sc_hd__nand3_4 _34909_ (.A(_12547_),
    .B(_12553_),
    .C(_12556_),
    .Y(_12557_));
 sky130_fd_sc_hd__o21ai_2 _34910_ (.A1(_12202_),
    .A2(_12198_),
    .B1(_12204_),
    .Y(_12558_));
 sky130_fd_sc_hd__o21ai_2 _34911_ (.A1(_12554_),
    .A2(_12555_),
    .B1(_12551_),
    .Y(_12559_));
 sky130_fd_sc_hd__nand3_2 _34912_ (.A(_12549_),
    .B(_12550_),
    .C(_12552_),
    .Y(_12560_));
 sky130_fd_sc_hd__nand3_4 _34913_ (.A(_12558_),
    .B(_12559_),
    .C(_12560_),
    .Y(_12561_));
 sky130_fd_sc_hd__nor2_4 _34914_ (.A(_12048_),
    .B(_12046_),
    .Y(_12562_));
 sky130_fd_sc_hd__o2bb2ai_4 _34915_ (.A1_N(_12557_),
    .A2_N(_12561_),
    .B1(_12044_),
    .B2(_12562_),
    .Y(_12563_));
 sky130_fd_sc_hd__nor2_4 _34916_ (.A(_12044_),
    .B(_12562_),
    .Y(_12564_));
 sky130_fd_sc_hd__nand3_4 _34917_ (.A(_12557_),
    .B(_12561_),
    .C(_12564_),
    .Y(_12565_));
 sky130_fd_sc_hd__nand2_1 _34918_ (.A(_12053_),
    .B(_12058_),
    .Y(_12566_));
 sky130_fd_sc_hd__nand2_4 _34919_ (.A(_12566_),
    .B(_12057_),
    .Y(_12567_));
 sky130_fd_sc_hd__a21oi_4 _34920_ (.A1(_12563_),
    .A2(_12565_),
    .B1(_12567_),
    .Y(_12568_));
 sky130_fd_sc_hd__and3_1 _34921_ (.A(_12547_),
    .B(_12556_),
    .C(_12553_),
    .X(_12569_));
 sky130_fd_sc_hd__nand2_2 _34922_ (.A(_12561_),
    .B(_12564_),
    .Y(_12570_));
 sky130_fd_sc_hd__o211a_2 _34923_ (.A1(_12569_),
    .A2(_12570_),
    .B1(_12567_),
    .C1(_12563_),
    .X(_12571_));
 sky130_fd_sc_hd__o22ai_4 _34924_ (.A1(_12542_),
    .A2(_12546_),
    .B1(_12568_),
    .B2(_12571_),
    .Y(_12572_));
 sky130_fd_sc_hd__nand2_1 _34925_ (.A(_12214_),
    .B(_12223_),
    .Y(_12573_));
 sky130_fd_sc_hd__nand2_2 _34926_ (.A(_12573_),
    .B(_12218_),
    .Y(_12574_));
 sky130_fd_sc_hd__a21o_1 _34927_ (.A1(_12563_),
    .A2(_12565_),
    .B1(_12567_),
    .X(_12575_));
 sky130_fd_sc_hd__a21oi_4 _34928_ (.A1(_12526_),
    .A2(_12529_),
    .B1(_12530_),
    .Y(_12576_));
 sky130_fd_sc_hd__o21ai_1 _34929_ (.A1(_12576_),
    .A2(_12544_),
    .B1(_12541_),
    .Y(_12577_));
 sky130_fd_sc_hd__nand2_1 _34930_ (.A(_12536_),
    .B(_12539_),
    .Y(_12578_));
 sky130_fd_sc_hd__o21ai_1 _34931_ (.A1(_12533_),
    .A2(_12535_),
    .B1(_12537_),
    .Y(_12579_));
 sky130_fd_sc_hd__nand2_2 _34932_ (.A(_12578_),
    .B(_12579_),
    .Y(_12580_));
 sky130_fd_sc_hd__nand3_1 _34933_ (.A(_12531_),
    .B(_12532_),
    .C(_12580_),
    .Y(_12581_));
 sky130_fd_sc_hd__nand2_2 _34934_ (.A(_12577_),
    .B(_12581_),
    .Y(_12582_));
 sky130_fd_sc_hd__nand3_4 _34935_ (.A(_12563_),
    .B(_12567_),
    .C(_12565_),
    .Y(_12583_));
 sky130_fd_sc_hd__nand3_4 _34936_ (.A(_12575_),
    .B(_12582_),
    .C(_12583_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand3_4 _34937_ (.A(_12572_),
    .B(_12574_),
    .C(_12584_),
    .Y(_12585_));
 sky130_vsdinv _34938_ (.A(_12585_),
    .Y(_12586_));
 sky130_fd_sc_hd__o21a_1 _34939_ (.A1(_12104_),
    .A2(_12105_),
    .B1(_12065_),
    .X(_12587_));
 sky130_vsdinv _34940_ (.A(_12587_),
    .Y(_12588_));
 sky130_fd_sc_hd__o21ai_4 _34941_ (.A1(_12568_),
    .A2(_12571_),
    .B1(_12582_),
    .Y(_12589_));
 sky130_fd_sc_hd__a21boi_4 _34942_ (.A1(_12214_),
    .A2(_12223_),
    .B1_N(_12218_),
    .Y(_12590_));
 sky130_fd_sc_hd__o21ai_2 _34943_ (.A1(_12576_),
    .A2(_12544_),
    .B1(_12580_),
    .Y(_12591_));
 sky130_fd_sc_hd__o21ai_4 _34944_ (.A1(_12544_),
    .A2(_12545_),
    .B1(_12591_),
    .Y(_12592_));
 sky130_fd_sc_hd__nand3_4 _34945_ (.A(_12575_),
    .B(_12592_),
    .C(_12583_),
    .Y(_12593_));
 sky130_fd_sc_hd__nand3_4 _34946_ (.A(_12589_),
    .B(_12590_),
    .C(_12593_),
    .Y(_12594_));
 sky130_fd_sc_hd__nand2_2 _34947_ (.A(_12588_),
    .B(_12594_),
    .Y(_12595_));
 sky130_fd_sc_hd__nor2_2 _34948_ (.A(_12586_),
    .B(_12595_),
    .Y(_12596_));
 sky130_fd_sc_hd__nand2_1 _34949_ (.A(_12104_),
    .B(_12065_),
    .Y(_12597_));
 sky130_fd_sc_hd__a22oi_4 _34950_ (.A1(_12063_),
    .A2(_12597_),
    .B1(_12594_),
    .B2(_12585_),
    .Y(_12598_));
 sky130_fd_sc_hd__o2bb2ai_4 _34951_ (.A1_N(_12515_),
    .A2_N(_12522_),
    .B1(_12596_),
    .B2(_12598_),
    .Y(_12599_));
 sky130_fd_sc_hd__a31oi_4 _34952_ (.A1(_12589_),
    .A2(_12590_),
    .A3(_12593_),
    .B1(_12587_),
    .Y(_12600_));
 sky130_fd_sc_hd__a21oi_4 _34953_ (.A1(_12585_),
    .A2(_12600_),
    .B1(_12598_),
    .Y(_12601_));
 sky130_fd_sc_hd__nand3_4 _34954_ (.A(_12522_),
    .B(_12601_),
    .C(_12515_),
    .Y(_12602_));
 sky130_fd_sc_hd__nand3_4 _34955_ (.A(_12389_),
    .B(_12599_),
    .C(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__buf_2 _34956_ (.A(_12603_),
    .X(_12604_));
 sky130_fd_sc_hd__a2bb2oi_4 _34957_ (.A1_N(_12241_),
    .A2_N(_12388_),
    .B1(_12247_),
    .B2(_12243_),
    .Y(_12605_));
 sky130_fd_sc_hd__a21o_1 _34958_ (.A1(_12594_),
    .A2(_12585_),
    .B1(_12588_),
    .X(_12606_));
 sky130_fd_sc_hd__o21ai_2 _34959_ (.A1(_12586_),
    .A2(_12595_),
    .B1(_12606_),
    .Y(_12607_));
 sky130_fd_sc_hd__nand3_2 _34960_ (.A(_12522_),
    .B(_12515_),
    .C(_12607_),
    .Y(_12608_));
 sky130_fd_sc_hd__nand2_1 _34961_ (.A(_12522_),
    .B(_12515_),
    .Y(_12609_));
 sky130_fd_sc_hd__nand2_1 _34962_ (.A(_12609_),
    .B(_12601_),
    .Y(_12610_));
 sky130_fd_sc_hd__nand3_4 _34963_ (.A(_12605_),
    .B(_12608_),
    .C(_12610_),
    .Y(_12611_));
 sky130_vsdinv _34964_ (.A(_12268_),
    .Y(_12612_));
 sky130_fd_sc_hd__and2_1 _34965_ (.A(_12279_),
    .B(_12271_),
    .X(_12613_));
 sky130_fd_sc_hd__buf_8 _34966_ (.A(_11184_),
    .X(_12614_));
 sky130_fd_sc_hd__nand3_4 _34967_ (.A(_06447_),
    .B(_12614_),
    .C(net476),
    .Y(_12615_));
 sky130_fd_sc_hd__nand3_4 _34968_ (.A(_11186_),
    .B(_12614_),
    .C(_05780_),
    .Y(_12616_));
 sky130_vsdinv _34969_ (.A(_05772_),
    .Y(_12617_));
 sky130_vsdinv _34970_ (.A(\pcpi_mul.rs1[31] ),
    .Y(_12618_));
 sky130_fd_sc_hd__nor2_2 _34971_ (.A(_12617_),
    .B(_12618_),
    .Y(_12619_));
 sky130_fd_sc_hd__a21o_2 _34972_ (.A1(_12615_),
    .A2(_12616_),
    .B1(_12619_),
    .X(_12620_));
 sky130_fd_sc_hd__nand3_4 _34973_ (.A(_12619_),
    .B(_12615_),
    .C(_12616_),
    .Y(_12621_));
 sky130_fd_sc_hd__a21oi_4 _34974_ (.A1(_11189_),
    .A2(_12263_),
    .B1(_12262_),
    .Y(_12622_));
 sky130_fd_sc_hd__a21o_2 _34975_ (.A1(_12620_),
    .A2(_12621_),
    .B1(_12622_),
    .X(_12623_));
 sky130_fd_sc_hd__nand3_4 _34976_ (.A(_12620_),
    .B(_12622_),
    .C(_12621_),
    .Y(_12624_));
 sky130_fd_sc_hd__a21oi_2 _34977_ (.A1(_12623_),
    .A2(_12624_),
    .B1(_12282_),
    .Y(_12625_));
 sky130_fd_sc_hd__and3_1 _34978_ (.A(_12623_),
    .B(_12282_),
    .C(_12624_),
    .X(_12626_));
 sky130_fd_sc_hd__o22ai_4 _34979_ (.A1(_12612_),
    .A2(_12613_),
    .B1(_12625_),
    .B2(_12626_),
    .Y(_12627_));
 sky130_fd_sc_hd__a21o_1 _34980_ (.A1(_12623_),
    .A2(_12624_),
    .B1(_12282_),
    .X(_12628_));
 sky130_fd_sc_hd__nand2_1 _34981_ (.A(_12268_),
    .B(_12281_),
    .Y(_12629_));
 sky130_fd_sc_hd__nand2_1 _34982_ (.A(_12629_),
    .B(_12271_),
    .Y(_12630_));
 sky130_fd_sc_hd__nand3_4 _34983_ (.A(_12623_),
    .B(_12282_),
    .C(_12624_),
    .Y(_12631_));
 sky130_fd_sc_hd__nand3_4 _34984_ (.A(_12628_),
    .B(_12630_),
    .C(_12631_),
    .Y(_12632_));
 sky130_fd_sc_hd__a21oi_4 _34985_ (.A1(_12273_),
    .A2(_19677_),
    .B1(_11957_),
    .Y(_12633_));
 sky130_vsdinv _34986_ (.A(_12633_),
    .Y(_12634_));
 sky130_fd_sc_hd__clkbuf_4 _34987_ (.A(_12634_),
    .X(_12635_));
 sky130_fd_sc_hd__and3_1 _34988_ (.A(_12627_),
    .B(_12632_),
    .C(_12635_),
    .X(_12636_));
 sky130_fd_sc_hd__a21oi_4 _34989_ (.A1(_12627_),
    .A2(_12632_),
    .B1(_12635_),
    .Y(_12637_));
 sky130_fd_sc_hd__nor2_4 _34990_ (.A(_11205_),
    .B(_12295_),
    .Y(_12638_));
 sky130_fd_sc_hd__buf_4 _34991_ (.A(_09933_),
    .X(_12639_));
 sky130_fd_sc_hd__a22o_1 _34992_ (.A1(_05452_),
    .A2(_11179_),
    .B1(_05405_),
    .B2(_12639_),
    .X(_12640_));
 sky130_fd_sc_hd__nand2_2 _34993_ (.A(_19668_),
    .B(_11202_),
    .Y(_12641_));
 sky130_fd_sc_hd__nand3b_2 _34994_ (.A_N(_12638_),
    .B(_12640_),
    .C(_12641_),
    .Y(_12642_));
 sky130_fd_sc_hd__a21oi_2 _34995_ (.A1(_12084_),
    .A2(_12087_),
    .B1(_12082_),
    .Y(_12643_));
 sky130_fd_sc_hd__a22oi_4 _34996_ (.A1(_06493_),
    .A2(_10601_),
    .B1(_06505_),
    .B2(_12639_),
    .Y(_12644_));
 sky130_vsdinv _34997_ (.A(_12641_),
    .Y(_12645_));
 sky130_fd_sc_hd__o21ai_2 _34998_ (.A1(_12644_),
    .A2(_12638_),
    .B1(_12645_),
    .Y(_12646_));
 sky130_fd_sc_hd__nand3_4 _34999_ (.A(_12642_),
    .B(_12643_),
    .C(_12646_),
    .Y(_12647_));
 sky130_fd_sc_hd__nand3b_2 _35000_ (.A_N(_12638_),
    .B(_12640_),
    .C(_12645_),
    .Y(_12648_));
 sky130_fd_sc_hd__o22ai_4 _35001_ (.A1(_12080_),
    .A2(_12081_),
    .B1(_12083_),
    .B2(_12086_),
    .Y(_12649_));
 sky130_fd_sc_hd__o21ai_2 _35002_ (.A1(_12644_),
    .A2(_12638_),
    .B1(_12641_),
    .Y(_12650_));
 sky130_fd_sc_hd__nand3_4 _35003_ (.A(_12648_),
    .B(_12649_),
    .C(_12650_),
    .Y(_12651_));
 sky130_fd_sc_hd__nand2_1 _35004_ (.A(_12647_),
    .B(_12651_),
    .Y(_12652_));
 sky130_fd_sc_hd__a21oi_4 _35005_ (.A1(_12297_),
    .A2(_12302_),
    .B1(_12296_),
    .Y(_12653_));
 sky130_fd_sc_hd__nand2_4 _35006_ (.A(_12652_),
    .B(_12653_),
    .Y(_12654_));
 sky130_vsdinv _35007_ (.A(_12653_),
    .Y(_12655_));
 sky130_fd_sc_hd__nand3_4 _35008_ (.A(_12647_),
    .B(_12651_),
    .C(_12655_),
    .Y(_12656_));
 sky130_fd_sc_hd__nand2_1 _35009_ (.A(_12090_),
    .B(_12091_),
    .Y(_12657_));
 sky130_fd_sc_hd__nand2_2 _35010_ (.A(_12657_),
    .B(_12075_),
    .Y(_12658_));
 sky130_fd_sc_hd__a21oi_4 _35011_ (.A1(_12654_),
    .A2(_12656_),
    .B1(_12658_),
    .Y(_12659_));
 sky130_fd_sc_hd__and3_1 _35012_ (.A(_12066_),
    .B(_12072_),
    .C(_12074_),
    .X(_12660_));
 sky130_fd_sc_hd__o211a_1 _35013_ (.A1(_12660_),
    .A2(_12089_),
    .B1(_12656_),
    .C1(_12654_),
    .X(_12661_));
 sky130_fd_sc_hd__a21boi_4 _35014_ (.A1(_12304_),
    .A2(_12311_),
    .B1_N(_12308_),
    .Y(_12662_));
 sky130_fd_sc_hd__o21ai_4 _35015_ (.A1(_12659_),
    .A2(_12661_),
    .B1(_12662_),
    .Y(_12663_));
 sky130_fd_sc_hd__a21o_1 _35016_ (.A1(_12654_),
    .A2(_12656_),
    .B1(_12658_),
    .X(_12664_));
 sky130_fd_sc_hd__nand3_4 _35017_ (.A(_12654_),
    .B(_12658_),
    .C(_12656_),
    .Y(_12665_));
 sky130_fd_sc_hd__nand3b_4 _35018_ (.A_N(_12662_),
    .B(_12664_),
    .C(_12665_),
    .Y(_12666_));
 sky130_fd_sc_hd__o21ai_2 _35019_ (.A1(_12318_),
    .A2(_12313_),
    .B1(_12322_),
    .Y(_12667_));
 sky130_fd_sc_hd__a21oi_2 _35020_ (.A1(_12663_),
    .A2(_12666_),
    .B1(_12667_),
    .Y(_12668_));
 sky130_fd_sc_hd__nor2_1 _35021_ (.A(_12318_),
    .B(_12313_),
    .Y(_12669_));
 sky130_fd_sc_hd__o211a_1 _35022_ (.A1(_12316_),
    .A2(_12669_),
    .B1(_12666_),
    .C1(_12663_),
    .X(_12670_));
 sky130_fd_sc_hd__o22ai_4 _35023_ (.A1(_12636_),
    .A2(_12637_),
    .B1(_12668_),
    .B2(_12670_),
    .Y(_12671_));
 sky130_fd_sc_hd__nand2_1 _35024_ (.A(_12628_),
    .B(_12631_),
    .Y(_12672_));
 sky130_fd_sc_hd__and2_1 _35025_ (.A(_12629_),
    .B(_12271_),
    .X(_12673_));
 sky130_fd_sc_hd__a21oi_2 _35026_ (.A1(_12672_),
    .A2(_12673_),
    .B1(_12633_),
    .Y(_12674_));
 sky130_fd_sc_hd__a21oi_2 _35027_ (.A1(_12632_),
    .A2(_12674_),
    .B1(_12637_),
    .Y(_12675_));
 sky130_fd_sc_hd__nor2_1 _35028_ (.A(_12319_),
    .B(_12316_),
    .Y(_12676_));
 sky130_fd_sc_hd__o2bb2ai_2 _35029_ (.A1_N(_12666_),
    .A2_N(_12663_),
    .B1(_12313_),
    .B2(_12676_),
    .Y(_12677_));
 sky130_fd_sc_hd__nand3_4 _35030_ (.A(_12663_),
    .B(_12667_),
    .C(_12666_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand3_4 _35031_ (.A(_12675_),
    .B(_12677_),
    .C(_12678_),
    .Y(_12679_));
 sky130_fd_sc_hd__nand2_1 _35032_ (.A(_12671_),
    .B(_12679_),
    .Y(_12680_));
 sky130_fd_sc_hd__nor2_1 _35033_ (.A(_12098_),
    .B(_12246_),
    .Y(_12681_));
 sky130_fd_sc_hd__nand2_2 _35034_ (.A(_12680_),
    .B(_12681_),
    .Y(_12682_));
 sky130_fd_sc_hd__nand2_2 _35035_ (.A(_12110_),
    .B(_12113_),
    .Y(_12683_));
 sky130_fd_sc_hd__nand3_4 _35036_ (.A(_12683_),
    .B(_12671_),
    .C(_12679_),
    .Y(_12684_));
 sky130_fd_sc_hd__nand2_4 _35037_ (.A(_12338_),
    .B(_12328_),
    .Y(_12685_));
 sky130_fd_sc_hd__a21oi_1 _35038_ (.A1(_12682_),
    .A2(_12684_),
    .B1(_12685_),
    .Y(_12686_));
 sky130_fd_sc_hd__nand3_4 _35039_ (.A(_12682_),
    .B(_12685_),
    .C(_12684_),
    .Y(_12687_));
 sky130_vsdinv _35040_ (.A(_12687_),
    .Y(_12688_));
 sky130_fd_sc_hd__o2bb2ai_2 _35041_ (.A1_N(_12604_),
    .A2_N(_12611_),
    .B1(_12686_),
    .B2(_12688_),
    .Y(_12689_));
 sky130_fd_sc_hd__o211a_2 _35042_ (.A1(_12098_),
    .A2(_12246_),
    .B1(_12679_),
    .C1(_12671_),
    .X(_12690_));
 sky130_fd_sc_hd__nand2_4 _35043_ (.A(_12682_),
    .B(_12685_),
    .Y(_12691_));
 sky130_fd_sc_hd__a21oi_2 _35044_ (.A1(_12671_),
    .A2(_12679_),
    .B1(_12683_),
    .Y(_12692_));
 sky130_fd_sc_hd__o21bai_4 _35045_ (.A1(_12692_),
    .A2(_12690_),
    .B1_N(_12685_),
    .Y(_12693_));
 sky130_fd_sc_hd__o2111ai_4 _35046_ (.A1(_12690_),
    .A2(_12691_),
    .B1(_12693_),
    .C1(_12603_),
    .D1(_12611_),
    .Y(_12694_));
 sky130_vsdinv _35047_ (.A(_12249_),
    .Y(_12695_));
 sky130_fd_sc_hd__nand2_1 _35048_ (.A(_12238_),
    .B(_12239_),
    .Y(_12696_));
 sky130_fd_sc_hd__nand2_1 _35049_ (.A(_12336_),
    .B(_12339_),
    .Y(_12697_));
 sky130_fd_sc_hd__nand2_1 _35050_ (.A(_12697_),
    .B(_12341_),
    .Y(_12698_));
 sky130_fd_sc_hd__nand2_2 _35051_ (.A(_12698_),
    .B(_12344_),
    .Y(_12699_));
 sky130_fd_sc_hd__a21oi_4 _35052_ (.A1(_12238_),
    .A2(_12249_),
    .B1(_12239_),
    .Y(_12700_));
 sky130_fd_sc_hd__o22ai_4 _35053_ (.A1(_12695_),
    .A2(_12696_),
    .B1(_12699_),
    .B2(_12700_),
    .Y(_12701_));
 sky130_fd_sc_hd__a21oi_4 _35054_ (.A1(_12689_),
    .A2(_12694_),
    .B1(_12701_),
    .Y(_12702_));
 sky130_vsdinv _35055_ (.A(_12604_),
    .Y(_12703_));
 sky130_fd_sc_hd__nand3_1 _35056_ (.A(_12611_),
    .B(_12693_),
    .C(_12687_),
    .Y(_12704_));
 sky130_fd_sc_hd__o211a_1 _35057_ (.A1(_12703_),
    .A2(_12704_),
    .B1(_12689_),
    .C1(_12701_),
    .X(_12705_));
 sky130_fd_sc_hd__nand2_1 _35058_ (.A(_12292_),
    .B(_12284_),
    .Y(_12706_));
 sky130_vsdinv _35059_ (.A(_12706_),
    .Y(_12707_));
 sky130_vsdinv _35060_ (.A(_12339_),
    .Y(_12708_));
 sky130_fd_sc_hd__nor2_1 _35061_ (.A(_12708_),
    .B(_12349_),
    .Y(_12709_));
 sky130_fd_sc_hd__nor2_2 _35062_ (.A(_12707_),
    .B(_12709_),
    .Y(_12710_));
 sky130_fd_sc_hd__nand2_1 _35063_ (.A(_12709_),
    .B(_12707_),
    .Y(_12711_));
 sky130_fd_sc_hd__and2b_2 _35064_ (.A_N(_12710_),
    .B(_12711_),
    .X(_12712_));
 sky130_fd_sc_hd__o21ai_4 _35065_ (.A1(_12702_),
    .A2(_12705_),
    .B1(_12712_),
    .Y(_12713_));
 sky130_fd_sc_hd__nand2_1 _35066_ (.A(_12611_),
    .B(_12604_),
    .Y(_12714_));
 sky130_fd_sc_hd__nand2_2 _35067_ (.A(_12693_),
    .B(_12687_),
    .Y(_12715_));
 sky130_fd_sc_hd__nand2_1 _35068_ (.A(_12350_),
    .B(_12256_),
    .Y(_12716_));
 sky130_fd_sc_hd__a22oi_4 _35069_ (.A1(_12714_),
    .A2(_12715_),
    .B1(_12716_),
    .B2(_12250_),
    .Y(_12717_));
 sky130_fd_sc_hd__nand2_2 _35070_ (.A(_12717_),
    .B(_12694_),
    .Y(_12718_));
 sky130_fd_sc_hd__a22oi_4 _35071_ (.A1(_12693_),
    .A2(_12687_),
    .B1(_12611_),
    .B2(_12604_),
    .Y(_12719_));
 sky130_fd_sc_hd__o2111a_1 _35072_ (.A1(_12690_),
    .A2(_12691_),
    .B1(_12693_),
    .C1(_12604_),
    .D1(_12611_),
    .X(_12720_));
 sky130_fd_sc_hd__o21a_1 _35073_ (.A1(_12699_),
    .A2(_12700_),
    .B1(_12250_),
    .X(_12721_));
 sky130_fd_sc_hd__o21ai_4 _35074_ (.A1(_12719_),
    .A2(_12720_),
    .B1(_12721_),
    .Y(_12722_));
 sky130_vsdinv _35075_ (.A(_12710_),
    .Y(_12723_));
 sky130_fd_sc_hd__nand2_2 _35076_ (.A(_12723_),
    .B(_12711_),
    .Y(_12724_));
 sky130_fd_sc_hd__nand3_4 _35077_ (.A(_12718_),
    .B(_12722_),
    .C(_12724_),
    .Y(_12725_));
 sky130_fd_sc_hd__nand3_4 _35078_ (.A(_12387_),
    .B(_12713_),
    .C(_12725_),
    .Y(_12726_));
 sky130_fd_sc_hd__o21ai_2 _35079_ (.A1(_12702_),
    .A2(_12705_),
    .B1(_12724_),
    .Y(_12727_));
 sky130_fd_sc_hd__nand3_4 _35080_ (.A(_12718_),
    .B(_12722_),
    .C(_12712_),
    .Y(_12728_));
 sky130_fd_sc_hd__o21ai_2 _35081_ (.A1(_12367_),
    .A2(_12354_),
    .B1(_12366_),
    .Y(_12729_));
 sky130_fd_sc_hd__nand3_4 _35082_ (.A(_12727_),
    .B(_12728_),
    .C(_12729_),
    .Y(_12730_));
 sky130_fd_sc_hd__a21oi_1 _35083_ (.A1(_12726_),
    .A2(_12730_),
    .B1(_12370_),
    .Y(_12731_));
 sky130_fd_sc_hd__and3_1 _35084_ (.A(_12726_),
    .B(_12730_),
    .C(_12370_),
    .X(_12732_));
 sky130_fd_sc_hd__nand2_1 _35085_ (.A(_12369_),
    .B(_12022_),
    .Y(_12733_));
 sky130_fd_sc_hd__nand2_2 _35086_ (.A(_12733_),
    .B(_12374_),
    .Y(_12734_));
 sky130_fd_sc_hd__o21bai_2 _35087_ (.A1(_12731_),
    .A2(_12732_),
    .B1_N(_12734_),
    .Y(_12735_));
 sky130_fd_sc_hd__a21o_1 _35088_ (.A1(_12726_),
    .A2(_12730_),
    .B1(_12370_),
    .X(_12736_));
 sky130_fd_sc_hd__nand3_2 _35089_ (.A(_12726_),
    .B(_12730_),
    .C(_12370_),
    .Y(_12737_));
 sky130_fd_sc_hd__nand3_4 _35090_ (.A(_12736_),
    .B(_12734_),
    .C(_12737_),
    .Y(_12738_));
 sky130_fd_sc_hd__and2_1 _35091_ (.A(_12735_),
    .B(_12738_),
    .X(_12739_));
 sky130_vsdinv _35092_ (.A(_12739_),
    .Y(_12740_));
 sky130_fd_sc_hd__nand2_8 _35093_ (.A(_12040_),
    .B(_11677_),
    .Y(_12741_));
 sky130_fd_sc_hd__o2111ai_4 _35094_ (.A1(_12376_),
    .A2(_12380_),
    .B1(_12038_),
    .C1(_12034_),
    .D1(_12383_),
    .Y(_12742_));
 sky130_fd_sc_hd__a21oi_1 _35095_ (.A1(_12381_),
    .A2(_12375_),
    .B1(_12382_),
    .Y(_12743_));
 sky130_fd_sc_hd__o22ai_1 _35096_ (.A1(_12376_),
    .A2(_12380_),
    .B1(_12038_),
    .B2(_12743_),
    .Y(_12744_));
 sky130_fd_sc_hd__o21bai_4 _35097_ (.A1(_12741_),
    .A2(_12742_),
    .B1_N(_12744_),
    .Y(_12745_));
 sky130_fd_sc_hd__nand3_1 _35098_ (.A(_12041_),
    .B(_12039_),
    .C(_12384_),
    .Y(_12746_));
 sky130_fd_sc_hd__and2b_1 _35099_ (.A_N(_12746_),
    .B(net409),
    .X(_12747_));
 sky130_fd_sc_hd__nor2_2 _35100_ (.A(_12745_),
    .B(_12747_),
    .Y(_12748_));
 sky130_fd_sc_hd__or2_1 _35101_ (.A(_12740_),
    .B(_12748_),
    .X(_12749_));
 sky130_fd_sc_hd__nand2_1 _35102_ (.A(_12748_),
    .B(_12740_),
    .Y(_12750_));
 sky130_fd_sc_hd__and2_4 _35103_ (.A(_12749_),
    .B(_12750_),
    .X(_02655_));
 sky130_fd_sc_hd__nand2_1 _35104_ (.A(_12522_),
    .B(_12601_),
    .Y(_12751_));
 sky130_fd_sc_hd__nand2_2 _35105_ (.A(_12751_),
    .B(_12515_),
    .Y(_12752_));
 sky130_fd_sc_hd__nand3_4 _35106_ (.A(_11080_),
    .B(_10830_),
    .C(_05291_),
    .Y(_12753_));
 sky130_fd_sc_hd__nand2_1 _35107_ (.A(_10830_),
    .B(_05486_),
    .Y(_12754_));
 sky130_fd_sc_hd__o21ai_4 _35108_ (.A1(_19917_),
    .A2(_18474_),
    .B1(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__o21ai_4 _35109_ (.A1(_19918_),
    .A2(_12753_),
    .B1(_12755_),
    .Y(_12756_));
 sky130_fd_sc_hd__nand2_4 _35110_ (.A(net498),
    .B(_05481_),
    .Y(_12757_));
 sky130_vsdinv _35111_ (.A(_12757_),
    .Y(_12758_));
 sky130_fd_sc_hd__nand2_1 _35112_ (.A(_12756_),
    .B(_12758_),
    .Y(_12759_));
 sky130_fd_sc_hd__o21ai_1 _35113_ (.A1(_05237_),
    .A2(_12393_),
    .B1(_12397_),
    .Y(_12760_));
 sky130_fd_sc_hd__nand2_2 _35114_ (.A(_12760_),
    .B(_12395_),
    .Y(_12761_));
 sky130_fd_sc_hd__nor2_4 _35115_ (.A(_05493_),
    .B(_12753_),
    .Y(_12762_));
 sky130_fd_sc_hd__nand3b_2 _35116_ (.A_N(_12762_),
    .B(_12755_),
    .C(_12757_),
    .Y(_12763_));
 sky130_fd_sc_hd__nand3_4 _35117_ (.A(_12759_),
    .B(_12761_),
    .C(_12763_),
    .Y(_12764_));
 sky130_fd_sc_hd__nand2_2 _35118_ (.A(_11348_),
    .B(_06105_),
    .Y(_12765_));
 sky130_fd_sc_hd__nand2_2 _35119_ (.A(_10046_),
    .B(_05796_),
    .Y(_12766_));
 sky130_fd_sc_hd__nor2_4 _35120_ (.A(_12765_),
    .B(_12766_),
    .Y(_12767_));
 sky130_fd_sc_hd__and2_1 _35121_ (.A(_12765_),
    .B(_12766_),
    .X(_12768_));
 sky130_fd_sc_hd__nand2_2 _35122_ (.A(_19591_),
    .B(_19901_),
    .Y(_12769_));
 sky130_vsdinv _35123_ (.A(_12769_),
    .Y(_12770_));
 sky130_fd_sc_hd__o21ai_1 _35124_ (.A1(_12767_),
    .A2(_12768_),
    .B1(_12770_),
    .Y(_12771_));
 sky130_fd_sc_hd__or2_1 _35125_ (.A(_12765_),
    .B(_12766_),
    .X(_12772_));
 sky130_fd_sc_hd__nand2_2 _35126_ (.A(_12765_),
    .B(_12766_),
    .Y(_12773_));
 sky130_fd_sc_hd__nand3_2 _35127_ (.A(_12772_),
    .B(_12769_),
    .C(_12773_),
    .Y(_12774_));
 sky130_fd_sc_hd__nand2_2 _35128_ (.A(_12771_),
    .B(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__nand2_2 _35129_ (.A(_12764_),
    .B(_12775_),
    .Y(_12776_));
 sky130_fd_sc_hd__nand2_1 _35130_ (.A(_12756_),
    .B(_12757_),
    .Y(_12777_));
 sky130_fd_sc_hd__nand3b_4 _35131_ (.A_N(_12762_),
    .B(_12755_),
    .C(_12758_),
    .Y(_12778_));
 sky130_fd_sc_hd__buf_6 _35132_ (.A(_11079_),
    .X(_12779_));
 sky130_fd_sc_hd__buf_6 _35133_ (.A(_11075_),
    .X(_12780_));
 sky130_fd_sc_hd__buf_6 _35134_ (.A(_12780_),
    .X(_12781_));
 sky130_fd_sc_hd__a22oi_4 _35135_ (.A1(_12779_),
    .A2(_19918_),
    .B1(_07426_),
    .B2(_12781_),
    .Y(_12782_));
 sky130_fd_sc_hd__o22ai_4 _35136_ (.A1(_19921_),
    .A2(_12393_),
    .B1(_12397_),
    .B2(_12782_),
    .Y(_12783_));
 sky130_fd_sc_hd__nand3_4 _35137_ (.A(_12777_),
    .B(_12778_),
    .C(_12783_),
    .Y(_12784_));
 sky130_vsdinv _35138_ (.A(_12784_),
    .Y(_12785_));
 sky130_fd_sc_hd__nor2_1 _35139_ (.A(_12767_),
    .B(_12768_),
    .Y(_12786_));
 sky130_fd_sc_hd__nor2_1 _35140_ (.A(_12770_),
    .B(_12786_),
    .Y(_12787_));
 sky130_fd_sc_hd__nand2_1 _35141_ (.A(_12772_),
    .B(_12773_),
    .Y(_12788_));
 sky130_fd_sc_hd__nor2_1 _35142_ (.A(_12769_),
    .B(_12788_),
    .Y(_12789_));
 sky130_fd_sc_hd__o2bb2ai_2 _35143_ (.A1_N(_12784_),
    .A2_N(_12764_),
    .B1(_12787_),
    .B2(_12789_),
    .Y(_12790_));
 sky130_fd_sc_hd__nand2_1 _35144_ (.A(_12410_),
    .B(_12426_),
    .Y(_12791_));
 sky130_fd_sc_hd__nand2_1 _35145_ (.A(_12791_),
    .B(_12405_),
    .Y(_12792_));
 sky130_fd_sc_hd__o211ai_4 _35146_ (.A1(_12776_),
    .A2(_12785_),
    .B1(_12790_),
    .C1(_12792_),
    .Y(_12793_));
 sky130_vsdinv _35147_ (.A(_12771_),
    .Y(_12794_));
 sky130_vsdinv _35148_ (.A(_12774_),
    .Y(_12795_));
 sky130_fd_sc_hd__o2bb2ai_4 _35149_ (.A1_N(_12784_),
    .A2_N(_12764_),
    .B1(_12794_),
    .B2(_12795_),
    .Y(_12796_));
 sky130_fd_sc_hd__nand3b_4 _35150_ (.A_N(_12775_),
    .B(_12784_),
    .C(_12764_),
    .Y(_12797_));
 sky130_fd_sc_hd__a21oi_2 _35151_ (.A1(_12396_),
    .A2(_12397_),
    .B1(_12408_),
    .Y(_12798_));
 sky130_fd_sc_hd__a22oi_4 _35152_ (.A1(_12798_),
    .A2(_12400_),
    .B1(_12410_),
    .B2(_12426_),
    .Y(_12799_));
 sky130_fd_sc_hd__nand3_4 _35153_ (.A(_12796_),
    .B(_12797_),
    .C(_12799_),
    .Y(_12800_));
 sky130_fd_sc_hd__nand2_1 _35154_ (.A(_12793_),
    .B(_12800_),
    .Y(_12801_));
 sky130_fd_sc_hd__a22oi_4 _35155_ (.A1(_09485_),
    .A2(_05977_),
    .B1(_19600_),
    .B2(_06116_),
    .Y(_12802_));
 sky130_fd_sc_hd__nand3_4 _35156_ (.A(_10260_),
    .B(_10257_),
    .C(_06649_),
    .Y(_12803_));
 sky130_fd_sc_hd__nor2_8 _35157_ (.A(net443),
    .B(_12803_),
    .Y(_12804_));
 sky130_fd_sc_hd__nand2_2 _35158_ (.A(_11801_),
    .B(_06462_),
    .Y(_12805_));
 sky130_vsdinv _35159_ (.A(_12805_),
    .Y(_12806_));
 sky130_fd_sc_hd__o21ai_2 _35160_ (.A1(_12802_),
    .A2(_12804_),
    .B1(_12806_),
    .Y(_12807_));
 sky130_fd_sc_hd__a21oi_4 _35161_ (.A1(_12416_),
    .A2(_12420_),
    .B1(_12414_),
    .Y(_12808_));
 sky130_fd_sc_hd__a22o_1 _35162_ (.A1(_19597_),
    .A2(_06119_),
    .B1(_19600_),
    .B2(_06289_),
    .X(_12809_));
 sky130_fd_sc_hd__o211ai_2 _35163_ (.A1(_06471_),
    .A2(_12803_),
    .B1(_12805_),
    .C1(_12809_),
    .Y(_12810_));
 sky130_fd_sc_hd__nand3_4 _35164_ (.A(_12807_),
    .B(_12808_),
    .C(_12810_),
    .Y(_12811_));
 sky130_fd_sc_hd__o21ai_2 _35165_ (.A1(_12802_),
    .A2(_12804_),
    .B1(_12805_),
    .Y(_12812_));
 sky130_fd_sc_hd__o21ai_2 _35166_ (.A1(_12415_),
    .A2(_12411_),
    .B1(_12419_),
    .Y(_12813_));
 sky130_fd_sc_hd__o211ai_2 _35167_ (.A1(_06471_),
    .A2(_12803_),
    .B1(_12806_),
    .C1(_12809_),
    .Y(_12814_));
 sky130_fd_sc_hd__nand3_4 _35168_ (.A(_12812_),
    .B(_12813_),
    .C(_12814_),
    .Y(_12815_));
 sky130_fd_sc_hd__a21oi_2 _35169_ (.A1(_12440_),
    .A2(_12442_),
    .B1(_12439_),
    .Y(_12816_));
 sky130_vsdinv _35170_ (.A(_12816_),
    .Y(_12817_));
 sky130_fd_sc_hd__a21oi_4 _35171_ (.A1(_12811_),
    .A2(_12815_),
    .B1(_12817_),
    .Y(_12818_));
 sky130_fd_sc_hd__and3_2 _35172_ (.A(_12811_),
    .B(_12815_),
    .C(_12817_),
    .X(_12819_));
 sky130_fd_sc_hd__nor2_8 _35173_ (.A(_12818_),
    .B(_12819_),
    .Y(_12820_));
 sky130_fd_sc_hd__nand2_1 _35174_ (.A(_12801_),
    .B(_12820_),
    .Y(_12821_));
 sky130_fd_sc_hd__a21boi_4 _35175_ (.A1(_12428_),
    .A2(_12456_),
    .B1_N(_12436_),
    .Y(_12822_));
 sky130_fd_sc_hd__nand3b_2 _35176_ (.A_N(_12820_),
    .B(_12793_),
    .C(_12800_),
    .Y(_12823_));
 sky130_fd_sc_hd__nand3_4 _35177_ (.A(_12821_),
    .B(_12822_),
    .C(_12823_),
    .Y(_12824_));
 sky130_fd_sc_hd__nand2_1 _35178_ (.A(_12456_),
    .B(_12428_),
    .Y(_12825_));
 sky130_fd_sc_hd__nand2_4 _35179_ (.A(_12825_),
    .B(_12436_),
    .Y(_12826_));
 sky130_fd_sc_hd__o2bb2ai_4 _35180_ (.A1_N(_12800_),
    .A2_N(_12793_),
    .B1(_12818_),
    .B2(_12819_),
    .Y(_12827_));
 sky130_fd_sc_hd__nand3_4 _35181_ (.A(_12793_),
    .B(_12820_),
    .C(_12800_),
    .Y(_12828_));
 sky130_fd_sc_hd__nand3_4 _35182_ (.A(_12826_),
    .B(_12827_),
    .C(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__nand2_4 _35183_ (.A(_07757_),
    .B(_07343_),
    .Y(_12830_));
 sky130_fd_sc_hd__nand2_4 _35184_ (.A(_08567_),
    .B(_09607_),
    .Y(_12831_));
 sky130_fd_sc_hd__nor2_8 _35185_ (.A(_12830_),
    .B(_12831_),
    .Y(_12832_));
 sky130_fd_sc_hd__and2_2 _35186_ (.A(_12830_),
    .B(_12831_),
    .X(_12833_));
 sky130_fd_sc_hd__nand2_4 _35187_ (.A(_19627_),
    .B(_10394_),
    .Y(_12834_));
 sky130_fd_sc_hd__o21a_1 _35188_ (.A1(_12832_),
    .A2(_12833_),
    .B1(_12834_),
    .X(_12835_));
 sky130_fd_sc_hd__nor3_4 _35189_ (.A(_12834_),
    .B(_12832_),
    .C(_12833_),
    .Y(_12836_));
 sky130_fd_sc_hd__nand2_2 _35190_ (.A(_08549_),
    .B(_07642_),
    .Y(_12837_));
 sky130_fd_sc_hd__nand2_2 _35191_ (.A(_10066_),
    .B(_06634_),
    .Y(_12838_));
 sky130_fd_sc_hd__nor2_4 _35192_ (.A(_12837_),
    .B(_12838_),
    .Y(_12839_));
 sky130_fd_sc_hd__nand2_2 _35193_ (.A(_12837_),
    .B(_12838_),
    .Y(_12840_));
 sky130_fd_sc_hd__nand2_2 _35194_ (.A(_12470_),
    .B(_07052_),
    .Y(_12841_));
 sky130_vsdinv _35195_ (.A(_12841_),
    .Y(_12842_));
 sky130_fd_sc_hd__nand3b_2 _35196_ (.A_N(_12839_),
    .B(_12840_),
    .C(_12842_),
    .Y(_12843_));
 sky130_fd_sc_hd__a22oi_4 _35197_ (.A1(_19608_),
    .A2(_11848_),
    .B1(_12466_),
    .B2(_07060_),
    .Y(_12844_));
 sky130_fd_sc_hd__o21ai_2 _35198_ (.A1(_12844_),
    .A2(_12839_),
    .B1(_12841_),
    .Y(_12845_));
 sky130_fd_sc_hd__o21ai_2 _35199_ (.A1(_12471_),
    .A2(_12467_),
    .B1(_12476_),
    .Y(_12846_));
 sky130_fd_sc_hd__nand3_4 _35200_ (.A(_12843_),
    .B(_12845_),
    .C(_12846_),
    .Y(_12847_));
 sky130_fd_sc_hd__nand3b_2 _35201_ (.A_N(_12839_),
    .B(_12840_),
    .C(_12841_),
    .Y(_12848_));
 sky130_fd_sc_hd__a21oi_2 _35202_ (.A1(_12477_),
    .A2(_12472_),
    .B1(_12469_),
    .Y(_12849_));
 sky130_fd_sc_hd__o21ai_2 _35203_ (.A1(_12844_),
    .A2(_12839_),
    .B1(_12842_),
    .Y(_12850_));
 sky130_fd_sc_hd__nand3_4 _35204_ (.A(_12848_),
    .B(_12849_),
    .C(_12850_),
    .Y(_12851_));
 sky130_fd_sc_hd__a2bb2oi_4 _35205_ (.A1_N(_12835_),
    .A2_N(_12836_),
    .B1(_12847_),
    .B2(_12851_),
    .Y(_12852_));
 sky130_vsdinv _35206_ (.A(_12834_),
    .Y(_12853_));
 sky130_fd_sc_hd__nor3_4 _35207_ (.A(_12853_),
    .B(_12832_),
    .C(_12833_),
    .Y(_12854_));
 sky130_fd_sc_hd__o21a_1 _35208_ (.A1(_12832_),
    .A2(_12833_),
    .B1(_12853_),
    .X(_12855_));
 sky130_fd_sc_hd__o211a_1 _35209_ (.A1(_12854_),
    .A2(_12855_),
    .B1(_12847_),
    .C1(_12851_),
    .X(_12856_));
 sky130_fd_sc_hd__nand2_1 _35210_ (.A(_12450_),
    .B(_12451_),
    .Y(_12857_));
 sky130_fd_sc_hd__nand2_4 _35211_ (.A(_12857_),
    .B(_12446_),
    .Y(_12858_));
 sky130_fd_sc_hd__o21bai_4 _35212_ (.A1(_12852_),
    .A2(_12856_),
    .B1_N(_12858_),
    .Y(_12859_));
 sky130_fd_sc_hd__nand2_1 _35213_ (.A(_12851_),
    .B(_12847_),
    .Y(_12860_));
 sky130_fd_sc_hd__nor2_2 _35214_ (.A(_12854_),
    .B(_12855_),
    .Y(_12861_));
 sky130_fd_sc_hd__nand2_2 _35215_ (.A(_12860_),
    .B(_12861_),
    .Y(_12862_));
 sky130_fd_sc_hd__o211ai_4 _35216_ (.A1(_12854_),
    .A2(_12855_),
    .B1(_12847_),
    .C1(_12851_),
    .Y(_12863_));
 sky130_fd_sc_hd__nand3_4 _35217_ (.A(_12862_),
    .B(_12858_),
    .C(_12863_),
    .Y(_12864_));
 sky130_fd_sc_hd__nand2_1 _35218_ (.A(_12490_),
    .B(_12479_),
    .Y(_12865_));
 sky130_fd_sc_hd__nand2_4 _35219_ (.A(_12865_),
    .B(_12494_),
    .Y(_12866_));
 sky130_fd_sc_hd__a21oi_4 _35220_ (.A1(_12859_),
    .A2(_12864_),
    .B1(_12866_),
    .Y(_12867_));
 sky130_fd_sc_hd__nand2_1 _35221_ (.A(_12862_),
    .B(_12858_),
    .Y(_12868_));
 sky130_fd_sc_hd__o211a_1 _35222_ (.A1(_12856_),
    .A2(_12868_),
    .B1(_12866_),
    .C1(_12859_),
    .X(_12869_));
 sky130_fd_sc_hd__o2bb2ai_2 _35223_ (.A1_N(_12824_),
    .A2_N(_12829_),
    .B1(_12867_),
    .B2(_12869_),
    .Y(_12870_));
 sky130_vsdinv _35224_ (.A(_12457_),
    .Y(_12871_));
 sky130_fd_sc_hd__nand2_1 _35225_ (.A(_12392_),
    .B(_12454_),
    .Y(_12872_));
 sky130_fd_sc_hd__a21oi_2 _35226_ (.A1(_12454_),
    .A2(_12457_),
    .B1(_12392_),
    .Y(_12873_));
 sky130_fd_sc_hd__o22ai_4 _35227_ (.A1(_12871_),
    .A2(_12872_),
    .B1(_12520_),
    .B2(_12873_),
    .Y(_12874_));
 sky130_fd_sc_hd__nor2_4 _35228_ (.A(_12867_),
    .B(_12869_),
    .Y(_12875_));
 sky130_fd_sc_hd__nand3_4 _35229_ (.A(_12875_),
    .B(_12824_),
    .C(_12829_),
    .Y(_12876_));
 sky130_fd_sc_hd__nand3_4 _35230_ (.A(_12870_),
    .B(_12874_),
    .C(_12876_),
    .Y(_12877_));
 sky130_fd_sc_hd__nand2_1 _35231_ (.A(_12824_),
    .B(_12829_),
    .Y(_12878_));
 sky130_fd_sc_hd__nand2_1 _35232_ (.A(_12878_),
    .B(_12875_),
    .Y(_12879_));
 sky130_fd_sc_hd__a22oi_4 _35233_ (.A1(_12459_),
    .A2(_12463_),
    .B1(_12153_),
    .B2(_12391_),
    .Y(_12880_));
 sky130_fd_sc_hd__a22oi_4 _35234_ (.A1(_12880_),
    .A2(_12457_),
    .B1(_12513_),
    .B2(_12465_),
    .Y(_12881_));
 sky130_fd_sc_hd__a21o_1 _35235_ (.A1(_12859_),
    .A2(_12864_),
    .B1(_12866_),
    .X(_12882_));
 sky130_fd_sc_hd__nand3_1 _35236_ (.A(_12859_),
    .B(_12864_),
    .C(_12866_),
    .Y(_12883_));
 sky130_fd_sc_hd__nand2_1 _35237_ (.A(_12882_),
    .B(_12883_),
    .Y(_12884_));
 sky130_fd_sc_hd__nand3_2 _35238_ (.A(_12884_),
    .B(_12824_),
    .C(_12829_),
    .Y(_12885_));
 sky130_fd_sc_hd__nand3_4 _35239_ (.A(_12879_),
    .B(_12881_),
    .C(_12885_),
    .Y(_12886_));
 sky130_fd_sc_hd__a21oi_4 _35240_ (.A1(_12503_),
    .A2(_12504_),
    .B1(_12499_),
    .Y(_12887_));
 sky130_fd_sc_hd__a21o_1 _35241_ (.A1(_12528_),
    .A2(_12524_),
    .B1(_12527_),
    .X(_12888_));
 sky130_fd_sc_hd__and4_4 _35242_ (.A(_06606_),
    .B(_06898_),
    .C(_19854_),
    .D(_10453_),
    .X(_12889_));
 sky130_fd_sc_hd__a22o_2 _35243_ (.A1(_06342_),
    .A2(_09082_),
    .B1(_06618_),
    .B2(_09365_),
    .X(_12890_));
 sky130_fd_sc_hd__nand2_2 _35244_ (.A(_06349_),
    .B(_09362_),
    .Y(_12891_));
 sky130_vsdinv _35245_ (.A(_12891_),
    .Y(_12892_));
 sky130_fd_sc_hd__nand3b_4 _35246_ (.A_N(_12889_),
    .B(_12890_),
    .C(_12892_),
    .Y(_12893_));
 sky130_fd_sc_hd__a22oi_4 _35247_ (.A1(net445),
    .A2(_19859_),
    .B1(_06423_),
    .B2(_19855_),
    .Y(_12894_));
 sky130_fd_sc_hd__o21ai_2 _35248_ (.A1(_12894_),
    .A2(_12889_),
    .B1(_12891_),
    .Y(_12895_));
 sky130_fd_sc_hd__nand3_4 _35249_ (.A(_12888_),
    .B(_12893_),
    .C(_12895_),
    .Y(_12896_));
 sky130_fd_sc_hd__nand3b_2 _35250_ (.A_N(_12889_),
    .B(_12890_),
    .C(_12891_),
    .Y(_12897_));
 sky130_fd_sc_hd__a21oi_2 _35251_ (.A1(_12528_),
    .A2(_12524_),
    .B1(_12527_),
    .Y(_12898_));
 sky130_fd_sc_hd__o21ai_2 _35252_ (.A1(_12894_),
    .A2(_12889_),
    .B1(_12892_),
    .Y(_12899_));
 sky130_fd_sc_hd__nand3_4 _35253_ (.A(_12897_),
    .B(_12898_),
    .C(_12899_),
    .Y(_12900_));
 sky130_fd_sc_hd__nand2_1 _35254_ (.A(_12896_),
    .B(_12900_),
    .Y(_12901_));
 sky130_fd_sc_hd__buf_6 _35255_ (.A(_09805_),
    .X(_12902_));
 sky130_fd_sc_hd__a22oi_4 _35256_ (.A1(_10737_),
    .A2(_09359_),
    .B1(_06336_),
    .B2(_11178_),
    .Y(_12903_));
 sky130_fd_sc_hd__nand2_2 _35257_ (.A(_06156_),
    .B(_11228_),
    .Y(_12904_));
 sky130_fd_sc_hd__nand2_2 _35258_ (.A(_05883_),
    .B(_09950_),
    .Y(_12905_));
 sky130_fd_sc_hd__nor2_4 _35259_ (.A(_12904_),
    .B(_12905_),
    .Y(_12906_));
 sky130_fd_sc_hd__nor2_1 _35260_ (.A(_12903_),
    .B(_12906_),
    .Y(_12907_));
 sky130_fd_sc_hd__o21ai_2 _35261_ (.A1(net450),
    .A2(_12902_),
    .B1(_12907_),
    .Y(_12908_));
 sky130_fd_sc_hd__nor2_4 _35262_ (.A(_05616_),
    .B(_09805_),
    .Y(_12909_));
 sky130_fd_sc_hd__o21ai_2 _35263_ (.A1(_12903_),
    .A2(_12906_),
    .B1(_12909_),
    .Y(_12910_));
 sky130_fd_sc_hd__nand2_4 _35264_ (.A(_12908_),
    .B(_12910_),
    .Y(_12911_));
 sky130_fd_sc_hd__and2_1 _35265_ (.A(_12901_),
    .B(_12911_),
    .X(_12912_));
 sky130_fd_sc_hd__nor2_2 _35266_ (.A(_12911_),
    .B(_12901_),
    .Y(_12913_));
 sky130_fd_sc_hd__nand2_1 _35267_ (.A(_12482_),
    .B(_12483_),
    .Y(_12914_));
 sky130_fd_sc_hd__a31o_1 _35268_ (.A1(_12914_),
    .A2(_11003_),
    .A3(_19875_),
    .B1(_12484_),
    .X(_12915_));
 sky130_fd_sc_hd__buf_6 _35269_ (.A(_09765_),
    .X(_12916_));
 sky130_fd_sc_hd__nand3_4 _35270_ (.A(_07744_),
    .B(_07928_),
    .C(_19868_),
    .Y(_12917_));
 sky130_fd_sc_hd__nand2_2 _35271_ (.A(_07435_),
    .B(_10458_),
    .Y(_12918_));
 sky130_vsdinv _35272_ (.A(_12918_),
    .Y(_12919_));
 sky130_fd_sc_hd__a22o_2 _35273_ (.A1(_10998_),
    .A2(_10149_),
    .B1(_10999_),
    .B2(_19866_),
    .X(_12920_));
 sky130_fd_sc_hd__o211ai_4 _35274_ (.A1(_12916_),
    .A2(_12917_),
    .B1(_12919_),
    .C1(_12920_),
    .Y(_12921_));
 sky130_fd_sc_hd__a22oi_4 _35275_ (.A1(_10990_),
    .A2(_19869_),
    .B1(_10991_),
    .B2(_10738_),
    .Y(_12922_));
 sky130_fd_sc_hd__nor2_4 _35276_ (.A(_09764_),
    .B(_12917_),
    .Y(_12923_));
 sky130_fd_sc_hd__o21ai_2 _35277_ (.A1(_12922_),
    .A2(_12923_),
    .B1(_12918_),
    .Y(_12924_));
 sky130_fd_sc_hd__nand3_4 _35278_ (.A(_12915_),
    .B(_12921_),
    .C(_12924_),
    .Y(_12925_));
 sky130_fd_sc_hd__nand3b_2 _35279_ (.A_N(_12923_),
    .B(_12920_),
    .C(_12918_),
    .Y(_12926_));
 sky130_fd_sc_hd__a21oi_2 _35280_ (.A1(_12486_),
    .A2(_12914_),
    .B1(_12484_),
    .Y(_12927_));
 sky130_fd_sc_hd__o21ai_2 _35281_ (.A1(_12922_),
    .A2(_12923_),
    .B1(_12919_),
    .Y(_12928_));
 sky130_fd_sc_hd__nand3_4 _35282_ (.A(_12926_),
    .B(_12927_),
    .C(_12928_),
    .Y(_12929_));
 sky130_fd_sc_hd__nor2_4 _35283_ (.A(_12551_),
    .B(_12555_),
    .Y(_12930_));
 sky130_fd_sc_hd__o2bb2ai_4 _35284_ (.A1_N(_12925_),
    .A2_N(_12929_),
    .B1(_12554_),
    .B2(_12930_),
    .Y(_12931_));
 sky130_fd_sc_hd__nor2_2 _35285_ (.A(_12554_),
    .B(_12930_),
    .Y(_12932_));
 sky130_fd_sc_hd__nand3_4 _35286_ (.A(_12925_),
    .B(_12929_),
    .C(_12932_),
    .Y(_12933_));
 sky130_fd_sc_hd__nand2_4 _35287_ (.A(_12570_),
    .B(_12557_),
    .Y(_12934_));
 sky130_fd_sc_hd__a21oi_4 _35288_ (.A1(_12931_),
    .A2(_12933_),
    .B1(_12934_),
    .Y(_12935_));
 sky130_fd_sc_hd__and3_1 _35289_ (.A(_12915_),
    .B(_12924_),
    .C(_12921_),
    .X(_12936_));
 sky130_fd_sc_hd__nand2_1 _35290_ (.A(_12929_),
    .B(_12932_),
    .Y(_12937_));
 sky130_fd_sc_hd__o211a_4 _35291_ (.A1(_12936_),
    .A2(_12937_),
    .B1(_12934_),
    .C1(_12931_),
    .X(_12938_));
 sky130_fd_sc_hd__o22ai_4 _35292_ (.A1(_12912_),
    .A2(_12913_),
    .B1(_12935_),
    .B2(_12938_),
    .Y(_12939_));
 sky130_fd_sc_hd__a21o_2 _35293_ (.A1(_12931_),
    .A2(_12933_),
    .B1(_12934_),
    .X(_12940_));
 sky130_fd_sc_hd__nand3_4 _35294_ (.A(_12931_),
    .B(_12934_),
    .C(_12933_),
    .Y(_12941_));
 sky130_fd_sc_hd__a21o_1 _35295_ (.A1(_12896_),
    .A2(_12900_),
    .B1(_12911_),
    .X(_12942_));
 sky130_fd_sc_hd__nand3_4 _35296_ (.A(_12911_),
    .B(_12896_),
    .C(_12900_),
    .Y(_12943_));
 sky130_fd_sc_hd__nand2_4 _35297_ (.A(_12942_),
    .B(_12943_),
    .Y(_12944_));
 sky130_fd_sc_hd__nand3_4 _35298_ (.A(_12940_),
    .B(_12941_),
    .C(_12944_),
    .Y(_12945_));
 sky130_fd_sc_hd__nand3_4 _35299_ (.A(_12887_),
    .B(_12939_),
    .C(_12945_),
    .Y(_12946_));
 sky130_fd_sc_hd__o21ai_4 _35300_ (.A1(_12935_),
    .A2(_12938_),
    .B1(_12944_),
    .Y(_12947_));
 sky130_fd_sc_hd__and2_1 _35301_ (.A(_12942_),
    .B(_12943_),
    .X(_12948_));
 sky130_fd_sc_hd__nand3_4 _35302_ (.A(_12948_),
    .B(_12940_),
    .C(_12941_),
    .Y(_12949_));
 sky130_fd_sc_hd__o21ai_4 _35303_ (.A1(_12510_),
    .A2(_12511_),
    .B1(_12507_),
    .Y(_12950_));
 sky130_fd_sc_hd__nand3_4 _35304_ (.A(_12947_),
    .B(_12949_),
    .C(_12950_),
    .Y(_12951_));
 sky130_fd_sc_hd__o21ai_4 _35305_ (.A1(_12568_),
    .A2(_12592_),
    .B1(_12583_),
    .Y(_12952_));
 sky130_fd_sc_hd__a21oi_4 _35306_ (.A1(_12946_),
    .A2(_12951_),
    .B1(_12952_),
    .Y(_12953_));
 sky130_fd_sc_hd__and3_1 _35307_ (.A(_12946_),
    .B(_12951_),
    .C(_12952_),
    .X(_12954_));
 sky130_fd_sc_hd__o2bb2ai_1 _35308_ (.A1_N(_12877_),
    .A2_N(_12886_),
    .B1(_12953_),
    .B2(_12954_),
    .Y(_12955_));
 sky130_fd_sc_hd__nor2_4 _35309_ (.A(_12953_),
    .B(_12954_),
    .Y(_12956_));
 sky130_fd_sc_hd__nand3_2 _35310_ (.A(_12956_),
    .B(_12886_),
    .C(_12877_),
    .Y(_12957_));
 sky130_fd_sc_hd__nand3_4 _35311_ (.A(_12752_),
    .B(_12955_),
    .C(_12957_),
    .Y(_12958_));
 sky130_fd_sc_hd__nand2_1 _35312_ (.A(_12886_),
    .B(_12877_),
    .Y(_12959_));
 sky130_fd_sc_hd__nand2_1 _35313_ (.A(_12959_),
    .B(_12956_),
    .Y(_12960_));
 sky130_fd_sc_hd__a22oi_4 _35314_ (.A1(_12236_),
    .A2(_12226_),
    .B1(_12516_),
    .B2(_12520_),
    .Y(_12961_));
 sky130_fd_sc_hd__a22oi_4 _35315_ (.A1(_12961_),
    .A2(_12514_),
    .B1(_12522_),
    .B2(_12601_),
    .Y(_12962_));
 sky130_fd_sc_hd__a21oi_4 _35316_ (.A1(_12939_),
    .A2(_12945_),
    .B1(_12887_),
    .Y(_12963_));
 sky130_fd_sc_hd__nand2_1 _35317_ (.A(_12946_),
    .B(_12952_),
    .Y(_12964_));
 sky130_fd_sc_hd__a21o_1 _35318_ (.A1(_12946_),
    .A2(_12951_),
    .B1(_12952_),
    .X(_12965_));
 sky130_fd_sc_hd__o21ai_2 _35319_ (.A1(_12963_),
    .A2(_12964_),
    .B1(_12965_),
    .Y(_12966_));
 sky130_fd_sc_hd__nand3_2 _35320_ (.A(_12966_),
    .B(_12886_),
    .C(_12877_),
    .Y(_12967_));
 sky130_fd_sc_hd__nand3_4 _35321_ (.A(_12960_),
    .B(_12962_),
    .C(_12967_),
    .Y(_12968_));
 sky130_fd_sc_hd__nand3_4 _35322_ (.A(_05440_),
    .B(_05404_),
    .C(\pcpi_mul.rs1[30] ),
    .Y(_12969_));
 sky130_fd_sc_hd__nor2_8 _35323_ (.A(_11205_),
    .B(_12969_),
    .Y(_12970_));
 sky130_fd_sc_hd__a22o_2 _35324_ (.A1(_05837_),
    .A2(_19834_),
    .B1(_19665_),
    .B2(_10504_),
    .X(_12971_));
 sky130_fd_sc_hd__nand2_2 _35325_ (.A(_19667_),
    .B(\pcpi_mul.rs1[31] ),
    .Y(_12972_));
 sky130_fd_sc_hd__nand3b_4 _35326_ (.A_N(_12970_),
    .B(_12971_),
    .C(_12972_),
    .Y(_12973_));
 sky130_fd_sc_hd__a22o_1 _35327_ (.A1(_06398_),
    .A2(_19851_),
    .B1(_06399_),
    .B2(_09820_),
    .X(_12974_));
 sky130_fd_sc_hd__a21oi_2 _35328_ (.A1(_12974_),
    .A2(_12539_),
    .B1(_12535_),
    .Y(_12975_));
 sky130_fd_sc_hd__a22oi_4 _35329_ (.A1(_06076_),
    .A2(_19834_),
    .B1(_06835_),
    .B2(_10504_),
    .Y(_12976_));
 sky130_vsdinv _35330_ (.A(_12972_),
    .Y(_12977_));
 sky130_fd_sc_hd__o21ai_2 _35331_ (.A1(_12976_),
    .A2(_12970_),
    .B1(_12977_),
    .Y(_12978_));
 sky130_fd_sc_hd__nand3_4 _35332_ (.A(_12973_),
    .B(_12975_),
    .C(_12978_),
    .Y(_12979_));
 sky130_fd_sc_hd__nor2_2 _35333_ (.A(_12537_),
    .B(_12533_),
    .Y(_12980_));
 sky130_fd_sc_hd__o211ai_4 _35334_ (.A1(_11206_),
    .A2(_12969_),
    .B1(_12977_),
    .C1(_12971_),
    .Y(_12981_));
 sky130_fd_sc_hd__o21ai_2 _35335_ (.A1(_12976_),
    .A2(_12970_),
    .B1(_12972_),
    .Y(_12982_));
 sky130_fd_sc_hd__o211ai_4 _35336_ (.A1(_12535_),
    .A2(_12980_),
    .B1(_12981_),
    .C1(_12982_),
    .Y(_12983_));
 sky130_fd_sc_hd__a21o_2 _35337_ (.A1(_12640_),
    .A2(_12645_),
    .B1(_12638_),
    .X(_12984_));
 sky130_fd_sc_hd__a21oi_4 _35338_ (.A1(_12979_),
    .A2(_12983_),
    .B1(_12984_),
    .Y(_12985_));
 sky130_fd_sc_hd__and3_2 _35339_ (.A(_12979_),
    .B(_12983_),
    .C(_12984_),
    .X(_12986_));
 sky130_fd_sc_hd__a21oi_2 _35340_ (.A1(_12531_),
    .A2(_12541_),
    .B1(_12544_),
    .Y(_12987_));
 sky130_fd_sc_hd__o21ai_4 _35341_ (.A1(_12985_),
    .A2(_12986_),
    .B1(_12987_),
    .Y(_12988_));
 sky130_fd_sc_hd__o21ai_4 _35342_ (.A1(_12580_),
    .A2(_12576_),
    .B1(_12532_),
    .Y(_12989_));
 sky130_fd_sc_hd__nand3_4 _35343_ (.A(_12979_),
    .B(_12983_),
    .C(_12984_),
    .Y(_12990_));
 sky130_fd_sc_hd__a21o_1 _35344_ (.A1(_12979_),
    .A2(_12983_),
    .B1(_12984_),
    .X(_12991_));
 sky130_fd_sc_hd__nand3_4 _35345_ (.A(_12989_),
    .B(_12990_),
    .C(_12991_),
    .Y(_12992_));
 sky130_fd_sc_hd__nand2_2 _35346_ (.A(_12988_),
    .B(_12992_),
    .Y(_12993_));
 sky130_fd_sc_hd__a21boi_4 _35347_ (.A1(_12647_),
    .A2(_12655_),
    .B1_N(_12651_),
    .Y(_12994_));
 sky130_fd_sc_hd__nand2_8 _35348_ (.A(_12993_),
    .B(_12994_),
    .Y(_12995_));
 sky130_vsdinv _35349_ (.A(_12994_),
    .Y(_12996_));
 sky130_fd_sc_hd__nand3_4 _35350_ (.A(_12988_),
    .B(_12992_),
    .C(_12996_),
    .Y(_12997_));
 sky130_fd_sc_hd__o21ai_4 _35351_ (.A1(_12662_),
    .A2(_12659_),
    .B1(_12665_),
    .Y(_12998_));
 sky130_fd_sc_hd__a21o_2 _35352_ (.A1(_12995_),
    .A2(_12997_),
    .B1(_12998_),
    .X(_12999_));
 sky130_fd_sc_hd__nand3_4 _35353_ (.A(_12995_),
    .B(_12998_),
    .C(_12997_),
    .Y(_13000_));
 sky130_fd_sc_hd__a21oi_2 _35354_ (.A1(_12620_),
    .A2(_12621_),
    .B1(_12622_),
    .Y(_13001_));
 sky130_fd_sc_hd__a21o_1 _35355_ (.A1(_12281_),
    .A2(_12624_),
    .B1(_13001_),
    .X(_13002_));
 sky130_fd_sc_hd__nor2_8 _35356_ (.A(_06258_),
    .B(net476),
    .Y(_13003_));
 sky130_fd_sc_hd__a21oi_4 _35357_ (.A1(_13003_),
    .A2(_12617_),
    .B1(_18469_),
    .Y(_13004_));
 sky130_vsdinv _35358_ (.A(_13004_),
    .Y(_13005_));
 sky130_fd_sc_hd__o21ai_2 _35359_ (.A1(_19674_),
    .A2(_19687_),
    .B1(net455),
    .Y(_13006_));
 sky130_fd_sc_hd__buf_6 _35360_ (.A(_12618_),
    .X(_13007_));
 sky130_fd_sc_hd__a21oi_4 _35361_ (.A1(_19674_),
    .A2(_19687_),
    .B1(_13007_),
    .Y(_13008_));
 sky130_fd_sc_hd__nor2_2 _35362_ (.A(_13006_),
    .B(_13008_),
    .Y(_13009_));
 sky130_fd_sc_hd__o21ai_2 _35363_ (.A1(_13005_),
    .A2(_13009_),
    .B1(_12281_),
    .Y(_13010_));
 sky130_fd_sc_hd__o2111ai_4 _35364_ (.A1(_13008_),
    .A2(_13006_),
    .B1(_12277_),
    .C1(_13004_),
    .D1(_12276_),
    .Y(_13011_));
 sky130_fd_sc_hd__nand2_1 _35365_ (.A(_13010_),
    .B(_13011_),
    .Y(_13012_));
 sky130_fd_sc_hd__nand2_2 _35366_ (.A(_13002_),
    .B(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__a21oi_2 _35367_ (.A1(_12624_),
    .A2(_12281_),
    .B1(_13001_),
    .Y(_13014_));
 sky130_fd_sc_hd__nand3_4 _35368_ (.A(_13014_),
    .B(_13011_),
    .C(_13010_),
    .Y(_13015_));
 sky130_fd_sc_hd__a21o_1 _35369_ (.A1(_13013_),
    .A2(_13015_),
    .B1(_12635_),
    .X(_13016_));
 sky130_fd_sc_hd__nand3_2 _35370_ (.A(_13013_),
    .B(_12635_),
    .C(_13015_),
    .Y(_13017_));
 sky130_fd_sc_hd__nand2_4 _35371_ (.A(_13016_),
    .B(_13017_),
    .Y(_13018_));
 sky130_fd_sc_hd__a21boi_4 _35372_ (.A1(_12999_),
    .A2(_13000_),
    .B1_N(_13018_),
    .Y(_13019_));
 sky130_fd_sc_hd__a21oi_4 _35373_ (.A1(_12995_),
    .A2(_12997_),
    .B1(_12998_),
    .Y(_13020_));
 sky130_fd_sc_hd__and3_2 _35374_ (.A(_12995_),
    .B(_12998_),
    .C(_12997_),
    .X(_13021_));
 sky130_fd_sc_hd__nor3_4 _35375_ (.A(_13018_),
    .B(_13020_),
    .C(_13021_),
    .Y(_13022_));
 sky130_fd_sc_hd__nand2_2 _35376_ (.A(_12595_),
    .B(_12585_),
    .Y(_13023_));
 sky130_fd_sc_hd__o21bai_2 _35377_ (.A1(_13019_),
    .A2(_13022_),
    .B1_N(_13023_),
    .Y(_13024_));
 sky130_fd_sc_hd__o21ai_2 _35378_ (.A1(_13020_),
    .A2(_13021_),
    .B1(_13018_),
    .Y(_13025_));
 sky130_fd_sc_hd__a31oi_4 _35379_ (.A1(_12995_),
    .A2(_12998_),
    .A3(_12997_),
    .B1(_13018_),
    .Y(_13026_));
 sky130_fd_sc_hd__nand2_4 _35380_ (.A(_13026_),
    .B(_12999_),
    .Y(_13027_));
 sky130_fd_sc_hd__nand3_4 _35381_ (.A(_13025_),
    .B(_13027_),
    .C(_13023_),
    .Y(_13028_));
 sky130_fd_sc_hd__nand2_2 _35382_ (.A(_12679_),
    .B(_12678_),
    .Y(_13029_));
 sky130_fd_sc_hd__a21oi_2 _35383_ (.A1(_13024_),
    .A2(_13028_),
    .B1(_13029_),
    .Y(_13030_));
 sky130_fd_sc_hd__and3_1 _35384_ (.A(_13024_),
    .B(_13028_),
    .C(_13029_),
    .X(_13031_));
 sky130_fd_sc_hd__o2bb2ai_4 _35385_ (.A1_N(_12958_),
    .A2_N(_12968_),
    .B1(_13030_),
    .B2(_13031_),
    .Y(_13032_));
 sky130_fd_sc_hd__o2bb2ai_2 _35386_ (.A1_N(_12999_),
    .A2_N(_13026_),
    .B1(_12586_),
    .B2(_12600_),
    .Y(_13033_));
 sky130_fd_sc_hd__nor2_4 _35387_ (.A(_13019_),
    .B(_13033_),
    .Y(_13034_));
 sky130_fd_sc_hd__nand2_2 _35388_ (.A(_13024_),
    .B(_13029_),
    .Y(_13035_));
 sky130_fd_sc_hd__a21oi_2 _35389_ (.A1(_13025_),
    .A2(_13027_),
    .B1(_13023_),
    .Y(_13036_));
 sky130_fd_sc_hd__o21bai_4 _35390_ (.A1(_13034_),
    .A2(_13036_),
    .B1_N(_13029_),
    .Y(_13037_));
 sky130_fd_sc_hd__o2111ai_4 _35391_ (.A1(_13034_),
    .A2(_13035_),
    .B1(_13037_),
    .C1(_12958_),
    .D1(_12968_),
    .Y(_13038_));
 sky130_vsdinv _35392_ (.A(_12602_),
    .Y(_13039_));
 sky130_fd_sc_hd__nand2_1 _35393_ (.A(_12389_),
    .B(_12599_),
    .Y(_13040_));
 sky130_fd_sc_hd__a21oi_4 _35394_ (.A1(_12599_),
    .A2(_12602_),
    .B1(_12389_),
    .Y(_13041_));
 sky130_fd_sc_hd__o22ai_4 _35395_ (.A1(_13039_),
    .A2(_13040_),
    .B1(_13041_),
    .B2(_12715_),
    .Y(_13042_));
 sky130_fd_sc_hd__a21oi_4 _35396_ (.A1(_13032_),
    .A2(_13038_),
    .B1(_13042_),
    .Y(_13043_));
 sky130_vsdinv _35397_ (.A(_12958_),
    .Y(_13044_));
 sky130_fd_sc_hd__nand3_2 _35398_ (.A(_13024_),
    .B(_13028_),
    .C(_13029_),
    .Y(_13045_));
 sky130_fd_sc_hd__nand3_4 _35399_ (.A(_12968_),
    .B(_13037_),
    .C(_13045_),
    .Y(_13046_));
 sky130_fd_sc_hd__o211a_2 _35400_ (.A1(_13044_),
    .A2(_13046_),
    .B1(_13032_),
    .C1(_13042_),
    .X(_13047_));
 sky130_vsdinv _35401_ (.A(_12674_),
    .Y(_13048_));
 sky130_fd_sc_hd__nand2_2 _35402_ (.A(_13048_),
    .B(_12632_),
    .Y(_13049_));
 sky130_fd_sc_hd__nand2_4 _35403_ (.A(_12691_),
    .B(_12684_),
    .Y(_13050_));
 sky130_fd_sc_hd__nor2_4 _35404_ (.A(_13049_),
    .B(_13050_),
    .Y(_13051_));
 sky130_vsdinv _35405_ (.A(_13049_),
    .Y(_13052_));
 sky130_fd_sc_hd__and2_1 _35406_ (.A(_12691_),
    .B(_12684_),
    .X(_13053_));
 sky130_fd_sc_hd__nor2_2 _35407_ (.A(_13052_),
    .B(_13053_),
    .Y(_13054_));
 sky130_fd_sc_hd__nor2_4 _35408_ (.A(_13051_),
    .B(_13054_),
    .Y(_13055_));
 sky130_fd_sc_hd__o21ai_2 _35409_ (.A1(_13043_),
    .A2(_13047_),
    .B1(_13055_),
    .Y(_13056_));
 sky130_fd_sc_hd__a22oi_4 _35410_ (.A1(_12694_),
    .A2(_12717_),
    .B1(_12722_),
    .B2(_12712_),
    .Y(_13057_));
 sky130_fd_sc_hd__nand2_1 _35411_ (.A(_13032_),
    .B(_13038_),
    .Y(_13058_));
 sky130_fd_sc_hd__o21a_1 _35412_ (.A1(_13041_),
    .A2(_12715_),
    .B1(_12604_),
    .X(_13059_));
 sky130_fd_sc_hd__nand2_4 _35413_ (.A(_13058_),
    .B(_13059_),
    .Y(_13060_));
 sky130_fd_sc_hd__nand3_4 _35414_ (.A(_13042_),
    .B(_13032_),
    .C(_13038_),
    .Y(_13061_));
 sky130_fd_sc_hd__xor2_4 _35415_ (.A(_13052_),
    .B(_13050_),
    .X(_13062_));
 sky130_fd_sc_hd__nand3_4 _35416_ (.A(_13060_),
    .B(_13061_),
    .C(_13062_),
    .Y(_13063_));
 sky130_fd_sc_hd__nand3_2 _35417_ (.A(_13056_),
    .B(_13057_),
    .C(_13063_),
    .Y(_13064_));
 sky130_fd_sc_hd__buf_2 _35418_ (.A(_13054_),
    .X(_13065_));
 sky130_fd_sc_hd__o22ai_4 _35419_ (.A1(_13065_),
    .A2(_13051_),
    .B1(_13043_),
    .B2(_13047_),
    .Y(_13066_));
 sky130_fd_sc_hd__o2bb2ai_2 _35420_ (.A1_N(_12694_),
    .A2_N(_12717_),
    .B1(_12724_),
    .B2(_12702_),
    .Y(_13067_));
 sky130_fd_sc_hd__nand3_4 _35421_ (.A(_13060_),
    .B(_13061_),
    .C(_13055_),
    .Y(_13068_));
 sky130_fd_sc_hd__nand3_4 _35422_ (.A(_13066_),
    .B(_13067_),
    .C(_13068_),
    .Y(_13069_));
 sky130_fd_sc_hd__a21oi_2 _35423_ (.A1(_13064_),
    .A2(_13069_),
    .B1(_12710_),
    .Y(_13070_));
 sky130_fd_sc_hd__and3_2 _35424_ (.A(_13064_),
    .B(_13069_),
    .C(_12710_),
    .X(_13071_));
 sky130_fd_sc_hd__and3_1 _35425_ (.A(_12727_),
    .B(_12729_),
    .C(_12728_),
    .X(_13072_));
 sky130_vsdinv _35426_ (.A(_12370_),
    .Y(_13073_));
 sky130_fd_sc_hd__a31oi_4 _35427_ (.A1(_12387_),
    .A2(_12713_),
    .A3(_12725_),
    .B1(_13073_),
    .Y(_13074_));
 sky130_fd_sc_hd__nor2_2 _35428_ (.A(_13072_),
    .B(_13074_),
    .Y(_13075_));
 sky130_fd_sc_hd__o21ai_4 _35429_ (.A1(_13070_),
    .A2(_13071_),
    .B1(_13075_),
    .Y(_13076_));
 sky130_fd_sc_hd__a31oi_4 _35430_ (.A1(_13056_),
    .A2(_13057_),
    .A3(_13063_),
    .B1(_12723_),
    .Y(_13077_));
 sky130_fd_sc_hd__nand2_1 _35431_ (.A(_13077_),
    .B(_13069_),
    .Y(_13078_));
 sky130_fd_sc_hd__nand2_1 _35432_ (.A(_13064_),
    .B(_13069_),
    .Y(_13079_));
 sky130_fd_sc_hd__nand2_1 _35433_ (.A(_13079_),
    .B(_12723_),
    .Y(_13080_));
 sky130_fd_sc_hd__o211ai_2 _35434_ (.A1(_13072_),
    .A2(_13074_),
    .B1(_13078_),
    .C1(_13080_),
    .Y(_13081_));
 sky130_fd_sc_hd__and2_2 _35435_ (.A(_13076_),
    .B(_13081_),
    .X(_13082_));
 sky130_fd_sc_hd__nand2_2 _35436_ (.A(_12749_),
    .B(_12738_),
    .Y(_13083_));
 sky130_fd_sc_hd__xor2_4 _35437_ (.A(_13082_),
    .B(_13083_),
    .X(_02656_));
 sky130_fd_sc_hd__a21oi_2 _35438_ (.A1(_13060_),
    .A2(_13055_),
    .B1(_13047_),
    .Y(_13084_));
 sky130_fd_sc_hd__nand2_1 _35439_ (.A(_13015_),
    .B(_12635_),
    .Y(_13085_));
 sky130_fd_sc_hd__nand2_4 _35440_ (.A(_13085_),
    .B(_13013_),
    .Y(_13086_));
 sky130_fd_sc_hd__nand2_4 _35441_ (.A(_13035_),
    .B(_13028_),
    .Y(_13087_));
 sky130_vsdinv _35442_ (.A(_13087_),
    .Y(_13088_));
 sky130_fd_sc_hd__nor2_2 _35443_ (.A(_13086_),
    .B(_13088_),
    .Y(_13089_));
 sky130_fd_sc_hd__inv_4 _35444_ (.A(_13086_),
    .Y(_13090_));
 sky130_fd_sc_hd__nor2_2 _35445_ (.A(_13090_),
    .B(_13087_),
    .Y(_13091_));
 sky130_fd_sc_hd__a21boi_4 _35446_ (.A1(_12956_),
    .A2(_12886_),
    .B1_N(_12877_),
    .Y(_13092_));
 sky130_fd_sc_hd__a21oi_4 _35447_ (.A1(_12827_),
    .A2(_12828_),
    .B1(_12826_),
    .Y(_13093_));
 sky130_fd_sc_hd__o21ai_2 _35448_ (.A1(_12884_),
    .A2(_13093_),
    .B1(_12829_),
    .Y(_13094_));
 sky130_fd_sc_hd__nand2_1 _35449_ (.A(_12820_),
    .B(_12800_),
    .Y(_13095_));
 sky130_fd_sc_hd__nand2_4 _35450_ (.A(_13095_),
    .B(_12793_),
    .Y(_13096_));
 sky130_fd_sc_hd__a22oi_4 _35451_ (.A1(_12779_),
    .A2(_05671_),
    .B1(net451),
    .B2(_11292_),
    .Y(_13097_));
 sky130_fd_sc_hd__nand2_8 _35452_ (.A(_11079_),
    .B(_08198_),
    .Y(_13098_));
 sky130_fd_sc_hd__buf_4 _35453_ (.A(_18474_),
    .X(_13099_));
 sky130_fd_sc_hd__nor3_4 _35454_ (.A(_19914_),
    .B(_13098_),
    .C(_13099_),
    .Y(_13100_));
 sky130_fd_sc_hd__nand2_4 _35455_ (.A(_10828_),
    .B(_06686_),
    .Y(_13101_));
 sky130_vsdinv _35456_ (.A(_13101_),
    .Y(_13102_));
 sky130_fd_sc_hd__o21ai_2 _35457_ (.A1(_13097_),
    .A2(_13100_),
    .B1(_13102_),
    .Y(_13103_));
 sky130_fd_sc_hd__a21oi_2 _35458_ (.A1(_12755_),
    .A2(_12758_),
    .B1(_12762_),
    .Y(_13104_));
 sky130_fd_sc_hd__nand2_4 _35459_ (.A(_05278_),
    .B(_12402_),
    .Y(_13105_));
 sky130_fd_sc_hd__nand2_4 _35460_ (.A(_13105_),
    .B(_13098_),
    .Y(_13106_));
 sky130_fd_sc_hd__buf_6 _35461_ (.A(_12780_),
    .X(_13107_));
 sky130_fd_sc_hd__nand3b_4 _35462_ (.A_N(_13098_),
    .B(_13107_),
    .C(_05279_),
    .Y(_13108_));
 sky130_fd_sc_hd__nand3_2 _35463_ (.A(_13106_),
    .B(_13108_),
    .C(_13101_),
    .Y(_13109_));
 sky130_fd_sc_hd__nand3_4 _35464_ (.A(_13103_),
    .B(_13104_),
    .C(_13109_),
    .Y(_13110_));
 sky130_fd_sc_hd__o21ai_2 _35465_ (.A1(_13097_),
    .A2(_13100_),
    .B1(_13101_),
    .Y(_13111_));
 sky130_fd_sc_hd__a21o_1 _35466_ (.A1(_12755_),
    .A2(_12758_),
    .B1(_12762_),
    .X(_13112_));
 sky130_fd_sc_hd__nand3_4 _35467_ (.A(_13106_),
    .B(_13108_),
    .C(_13102_),
    .Y(_13113_));
 sky130_fd_sc_hd__nand3_4 _35468_ (.A(_13111_),
    .B(_13112_),
    .C(_13113_),
    .Y(_13114_));
 sky130_fd_sc_hd__a22oi_4 _35469_ (.A1(_11348_),
    .A2(_19904_),
    .B1(net494),
    .B2(_19901_),
    .Y(_13115_));
 sky130_fd_sc_hd__nand3_2 _35470_ (.A(_10281_),
    .B(_19587_),
    .C(_06257_),
    .Y(_13116_));
 sky130_fd_sc_hd__nor2_4 _35471_ (.A(net442),
    .B(_13116_),
    .Y(_13117_));
 sky130_fd_sc_hd__clkbuf_2 _35472_ (.A(_10044_),
    .X(_13118_));
 sky130_fd_sc_hd__nor2_4 _35473_ (.A(_13118_),
    .B(_07102_),
    .Y(_13119_));
 sky130_fd_sc_hd__o21ai_1 _35474_ (.A1(_13115_),
    .A2(_13117_),
    .B1(_13119_),
    .Y(_13120_));
 sky130_vsdinv _35475_ (.A(_13120_),
    .Y(_13121_));
 sky130_fd_sc_hd__a211o_1 _35476_ (.A1(_19593_),
    .A2(_19899_),
    .B1(_13115_),
    .C1(_13117_),
    .X(_13122_));
 sky130_vsdinv _35477_ (.A(_13122_),
    .Y(_13123_));
 sky130_fd_sc_hd__o2bb2ai_2 _35478_ (.A1_N(_13110_),
    .A2_N(_13114_),
    .B1(_13121_),
    .B2(_13123_),
    .Y(_13124_));
 sky130_fd_sc_hd__a21oi_4 _35479_ (.A1(_12756_),
    .A2(_12757_),
    .B1(_12761_),
    .Y(_13125_));
 sky130_fd_sc_hd__a22oi_4 _35480_ (.A1(_13125_),
    .A2(_12778_),
    .B1(_12764_),
    .B2(_12775_),
    .Y(_13126_));
 sky130_vsdinv _35481_ (.A(_13119_),
    .Y(_13127_));
 sky130_fd_sc_hd__o21ai_1 _35482_ (.A1(_13115_),
    .A2(_13117_),
    .B1(_13127_),
    .Y(_13128_));
 sky130_vsdinv _35483_ (.A(_13115_),
    .Y(_13129_));
 sky130_fd_sc_hd__nand3b_1 _35484_ (.A_N(_13117_),
    .B(_13129_),
    .C(_13119_),
    .Y(_13130_));
 sky130_fd_sc_hd__nand2_1 _35485_ (.A(_13128_),
    .B(_13130_),
    .Y(_13131_));
 sky130_fd_sc_hd__nand3_2 _35486_ (.A(_13114_),
    .B(_13110_),
    .C(_13131_),
    .Y(_13132_));
 sky130_fd_sc_hd__nand3_4 _35487_ (.A(_13124_),
    .B(_13126_),
    .C(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__nand2_1 _35488_ (.A(_13114_),
    .B(_13110_),
    .Y(_13134_));
 sky130_fd_sc_hd__nand2_1 _35489_ (.A(_13134_),
    .B(_13131_),
    .Y(_13135_));
 sky130_fd_sc_hd__nand2_1 _35490_ (.A(_12776_),
    .B(_12784_),
    .Y(_13136_));
 sky130_fd_sc_hd__nand2_2 _35491_ (.A(_13122_),
    .B(_13120_),
    .Y(_13137_));
 sky130_fd_sc_hd__nand3_2 _35492_ (.A(_13114_),
    .B(_13137_),
    .C(_13110_),
    .Y(_13138_));
 sky130_fd_sc_hd__nand3_4 _35493_ (.A(_13135_),
    .B(_13136_),
    .C(_13138_),
    .Y(_13139_));
 sky130_fd_sc_hd__o21ai_4 _35494_ (.A1(_12770_),
    .A2(_12767_),
    .B1(_12773_),
    .Y(_13140_));
 sky130_fd_sc_hd__nand2_4 _35495_ (.A(_19596_),
    .B(_07502_),
    .Y(_13141_));
 sky130_fd_sc_hd__nand2_4 _35496_ (.A(_09227_),
    .B(_06465_),
    .Y(_13142_));
 sky130_fd_sc_hd__nor2_4 _35497_ (.A(_13141_),
    .B(_13142_),
    .Y(_13143_));
 sky130_fd_sc_hd__and2_1 _35498_ (.A(_13141_),
    .B(_13142_),
    .X(_13144_));
 sky130_fd_sc_hd__nand2_2 _35499_ (.A(_11801_),
    .B(_07064_),
    .Y(_13145_));
 sky130_fd_sc_hd__o21ai_2 _35500_ (.A1(_13143_),
    .A2(_13144_),
    .B1(_13145_),
    .Y(_13146_));
 sky130_fd_sc_hd__nand2_2 _35501_ (.A(_13141_),
    .B(_13142_),
    .Y(_13147_));
 sky130_vsdinv _35502_ (.A(_13145_),
    .Y(_13148_));
 sky130_fd_sc_hd__nand3b_4 _35503_ (.A_N(_13143_),
    .B(_13147_),
    .C(_13148_),
    .Y(_13149_));
 sky130_fd_sc_hd__nand3b_4 _35504_ (.A_N(_13140_),
    .B(_13146_),
    .C(_13149_),
    .Y(_13150_));
 sky130_fd_sc_hd__o21ai_2 _35505_ (.A1(_13143_),
    .A2(_13144_),
    .B1(_13148_),
    .Y(_13151_));
 sky130_fd_sc_hd__nand3b_2 _35506_ (.A_N(_13143_),
    .B(_13147_),
    .C(_13145_),
    .Y(_13152_));
 sky130_fd_sc_hd__nand3_4 _35507_ (.A(_13151_),
    .B(_13152_),
    .C(_13140_),
    .Y(_13153_));
 sky130_fd_sc_hd__nor2_4 _35508_ (.A(_12805_),
    .B(_12802_),
    .Y(_13154_));
 sky130_fd_sc_hd__or2_2 _35509_ (.A(_12804_),
    .B(_13154_),
    .X(_13155_));
 sky130_fd_sc_hd__a21oi_4 _35510_ (.A1(_13150_),
    .A2(_13153_),
    .B1(_13155_),
    .Y(_13156_));
 sky130_fd_sc_hd__and3_2 _35511_ (.A(_13150_),
    .B(_13153_),
    .C(_13155_),
    .X(_13157_));
 sky130_fd_sc_hd__o2bb2ai_4 _35512_ (.A1_N(_13133_),
    .A2_N(_13139_),
    .B1(_13156_),
    .B2(_13157_),
    .Y(_13158_));
 sky130_fd_sc_hd__o21a_1 _35513_ (.A1(_12804_),
    .A2(_13154_),
    .B1(_13153_),
    .X(_13159_));
 sky130_fd_sc_hd__a21oi_4 _35514_ (.A1(_13159_),
    .A2(_13150_),
    .B1(_13156_),
    .Y(_13160_));
 sky130_fd_sc_hd__nand3_4 _35515_ (.A(_13160_),
    .B(_13139_),
    .C(_13133_),
    .Y(_13161_));
 sky130_fd_sc_hd__nand3_4 _35516_ (.A(_13096_),
    .B(_13158_),
    .C(_13161_),
    .Y(_13162_));
 sky130_fd_sc_hd__nand2_1 _35517_ (.A(_13139_),
    .B(_13133_),
    .Y(_13163_));
 sky130_fd_sc_hd__nand2_1 _35518_ (.A(_13163_),
    .B(_13160_),
    .Y(_13164_));
 sky130_fd_sc_hd__a21oi_4 _35519_ (.A1(_12796_),
    .A2(_12797_),
    .B1(_12799_),
    .Y(_13165_));
 sky130_fd_sc_hd__a21oi_4 _35520_ (.A1(_12820_),
    .A2(_12800_),
    .B1(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__o211ai_4 _35521_ (.A1(_13156_),
    .A2(_13157_),
    .B1(_13133_),
    .C1(_13139_),
    .Y(_13167_));
 sky130_fd_sc_hd__nand3_4 _35522_ (.A(_13164_),
    .B(_13166_),
    .C(_13167_),
    .Y(_13168_));
 sky130_fd_sc_hd__nand2_2 _35523_ (.A(_12861_),
    .B(_12847_),
    .Y(_13169_));
 sky130_fd_sc_hd__nand2_4 _35524_ (.A(_19607_),
    .B(_06443_),
    .Y(_13170_));
 sky130_fd_sc_hd__nand2_4 _35525_ (.A(_09680_),
    .B(_06654_),
    .Y(_13171_));
 sky130_fd_sc_hd__nor2_8 _35526_ (.A(_13170_),
    .B(_13171_),
    .Y(_13172_));
 sky130_fd_sc_hd__and2_1 _35527_ (.A(_13170_),
    .B(_13171_),
    .X(_13173_));
 sky130_fd_sc_hd__nand2_2 _35528_ (.A(_19616_),
    .B(_19877_),
    .Y(_13174_));
 sky130_fd_sc_hd__o21ai_2 _35529_ (.A1(_13172_),
    .A2(_13173_),
    .B1(_13174_),
    .Y(_13175_));
 sky130_fd_sc_hd__nand2_4 _35530_ (.A(_13170_),
    .B(_13171_),
    .Y(_13176_));
 sky130_vsdinv _35531_ (.A(_13174_),
    .Y(_13177_));
 sky130_fd_sc_hd__nand3b_2 _35532_ (.A_N(_13172_),
    .B(_13176_),
    .C(_13177_),
    .Y(_13178_));
 sky130_fd_sc_hd__a21o_1 _35533_ (.A1(_12842_),
    .A2(_12840_),
    .B1(_12839_),
    .X(_13179_));
 sky130_fd_sc_hd__nand3_4 _35534_ (.A(_13175_),
    .B(_13178_),
    .C(_13179_),
    .Y(_13180_));
 sky130_fd_sc_hd__o21ai_2 _35535_ (.A1(_13172_),
    .A2(_13173_),
    .B1(_13177_),
    .Y(_13181_));
 sky130_fd_sc_hd__nand3b_2 _35536_ (.A_N(_13172_),
    .B(_13176_),
    .C(_13174_),
    .Y(_13182_));
 sky130_fd_sc_hd__a21oi_2 _35537_ (.A1(_12842_),
    .A2(_12840_),
    .B1(_12839_),
    .Y(_13183_));
 sky130_fd_sc_hd__nand3_4 _35538_ (.A(_13181_),
    .B(_13182_),
    .C(_13183_),
    .Y(_13184_));
 sky130_fd_sc_hd__nand2_1 _35539_ (.A(_13180_),
    .B(_13184_),
    .Y(_13185_));
 sky130_fd_sc_hd__nand2_2 _35540_ (.A(_07934_),
    .B(_08735_),
    .Y(_13186_));
 sky130_fd_sc_hd__nand2_2 _35541_ (.A(_07758_),
    .B(_10394_),
    .Y(_13187_));
 sky130_fd_sc_hd__or2_2 _35542_ (.A(_13186_),
    .B(_13187_),
    .X(_13188_));
 sky130_fd_sc_hd__nand2_4 _35543_ (.A(_13186_),
    .B(_13187_),
    .Y(_13189_));
 sky130_fd_sc_hd__nand2_2 _35544_ (.A(_19628_),
    .B(_11724_),
    .Y(_13190_));
 sky130_fd_sc_hd__a21oi_2 _35545_ (.A1(_13188_),
    .A2(_13189_),
    .B1(_13190_),
    .Y(_13191_));
 sky130_fd_sc_hd__and3_1 _35546_ (.A(_13188_),
    .B(_13190_),
    .C(_13189_),
    .X(_13192_));
 sky130_fd_sc_hd__nor2_4 _35547_ (.A(_13191_),
    .B(_13192_),
    .Y(_13193_));
 sky130_fd_sc_hd__nand2_4 _35548_ (.A(_13185_),
    .B(_13193_),
    .Y(_13194_));
 sky130_fd_sc_hd__a21o_1 _35549_ (.A1(_13188_),
    .A2(_13189_),
    .B1(_13190_),
    .X(_13195_));
 sky130_fd_sc_hd__nand3_1 _35550_ (.A(_13188_),
    .B(_13190_),
    .C(_13189_),
    .Y(_13196_));
 sky130_fd_sc_hd__nand2_2 _35551_ (.A(_13195_),
    .B(_13196_),
    .Y(_13197_));
 sky130_fd_sc_hd__nand3_4 _35552_ (.A(_13197_),
    .B(_13180_),
    .C(_13184_),
    .Y(_13198_));
 sky130_fd_sc_hd__a21bo_2 _35553_ (.A1(_12811_),
    .A2(_12817_),
    .B1_N(_12815_),
    .X(_13199_));
 sky130_fd_sc_hd__a21o_1 _35554_ (.A1(_13194_),
    .A2(_13198_),
    .B1(_13199_),
    .X(_13200_));
 sky130_fd_sc_hd__nand3_4 _35555_ (.A(_13199_),
    .B(_13194_),
    .C(_13198_),
    .Y(_13201_));
 sky130_fd_sc_hd__a22oi_4 _35556_ (.A1(_12851_),
    .A2(_13169_),
    .B1(_13200_),
    .B2(_13201_),
    .Y(_13202_));
 sky130_fd_sc_hd__a21oi_4 _35557_ (.A1(_13194_),
    .A2(_13198_),
    .B1(_13199_),
    .Y(_13203_));
 sky130_fd_sc_hd__nand2_4 _35558_ (.A(_13169_),
    .B(_12851_),
    .Y(_13204_));
 sky130_vsdinv _35559_ (.A(_13201_),
    .Y(_13205_));
 sky130_fd_sc_hd__nor3_4 _35560_ (.A(_13203_),
    .B(_13204_),
    .C(_13205_),
    .Y(_13206_));
 sky130_fd_sc_hd__o2bb2ai_2 _35561_ (.A1_N(_13162_),
    .A2_N(_13168_),
    .B1(_13202_),
    .B2(_13206_),
    .Y(_13207_));
 sky130_fd_sc_hd__nor2_2 _35562_ (.A(_13204_),
    .B(_13203_),
    .Y(_13208_));
 sky130_fd_sc_hd__a21oi_4 _35563_ (.A1(_13201_),
    .A2(_13208_),
    .B1(_13202_),
    .Y(_13209_));
 sky130_fd_sc_hd__nand3_4 _35564_ (.A(_13209_),
    .B(_13168_),
    .C(_13162_),
    .Y(_13210_));
 sky130_fd_sc_hd__nand3_4 _35565_ (.A(_13094_),
    .B(_13207_),
    .C(_13210_),
    .Y(_13211_));
 sky130_fd_sc_hd__nand2_1 _35566_ (.A(_13168_),
    .B(_13162_),
    .Y(_13212_));
 sky130_fd_sc_hd__nand2_1 _35567_ (.A(_13212_),
    .B(_13209_),
    .Y(_13213_));
 sky130_fd_sc_hd__a21boi_4 _35568_ (.A1(_12875_),
    .A2(_12824_),
    .B1_N(_12829_),
    .Y(_13214_));
 sky130_fd_sc_hd__o21ai_1 _35569_ (.A1(_13203_),
    .A2(_13205_),
    .B1(_13204_),
    .Y(_13215_));
 sky130_fd_sc_hd__nand2_1 _35570_ (.A(_13208_),
    .B(_13201_),
    .Y(_13216_));
 sky130_fd_sc_hd__nand2_2 _35571_ (.A(_13215_),
    .B(_13216_),
    .Y(_13217_));
 sky130_fd_sc_hd__nand3_2 _35572_ (.A(_13217_),
    .B(_13168_),
    .C(_13162_),
    .Y(_13218_));
 sky130_fd_sc_hd__nand3_4 _35573_ (.A(_13213_),
    .B(_13214_),
    .C(_13218_),
    .Y(_13219_));
 sky130_fd_sc_hd__a21boi_4 _35574_ (.A1(_12859_),
    .A2(_12866_),
    .B1_N(_12864_),
    .Y(_13220_));
 sky130_fd_sc_hd__nand2_1 _35575_ (.A(_12830_),
    .B(_12831_),
    .Y(_13221_));
 sky130_fd_sc_hd__a21oi_4 _35576_ (.A1(_12853_),
    .A2(_13221_),
    .B1(_12832_),
    .Y(_13222_));
 sky130_fd_sc_hd__nand2_4 _35577_ (.A(_08615_),
    .B(_09772_),
    .Y(_13223_));
 sky130_fd_sc_hd__nand2_4 _35578_ (.A(_08873_),
    .B(_08337_),
    .Y(_13224_));
 sky130_fd_sc_hd__nor2_8 _35579_ (.A(_13223_),
    .B(_13224_),
    .Y(_13225_));
 sky130_fd_sc_hd__and2_4 _35580_ (.A(_13223_),
    .B(_13224_),
    .X(_13226_));
 sky130_fd_sc_hd__nand2_4 _35581_ (.A(_07435_),
    .B(_09082_),
    .Y(_13227_));
 sky130_fd_sc_hd__o21ai_2 _35582_ (.A1(_13225_),
    .A2(_13226_),
    .B1(_13227_),
    .Y(_13228_));
 sky130_fd_sc_hd__or2_2 _35583_ (.A(_13223_),
    .B(_13224_),
    .X(_13229_));
 sky130_fd_sc_hd__nand2_2 _35584_ (.A(_13223_),
    .B(_13224_),
    .Y(_13230_));
 sky130_vsdinv _35585_ (.A(_13227_),
    .Y(_13231_));
 sky130_fd_sc_hd__nand3_2 _35586_ (.A(_13229_),
    .B(_13230_),
    .C(_13231_),
    .Y(_13232_));
 sky130_fd_sc_hd__nand3b_4 _35587_ (.A_N(_13222_),
    .B(_13228_),
    .C(_13232_),
    .Y(_13233_));
 sky130_fd_sc_hd__o21ai_4 _35588_ (.A1(_13225_),
    .A2(_13226_),
    .B1(_13231_),
    .Y(_13234_));
 sky130_fd_sc_hd__nand3_4 _35589_ (.A(_13229_),
    .B(_13230_),
    .C(_13227_),
    .Y(_13235_));
 sky130_fd_sc_hd__nand3_1 _35590_ (.A(_13234_),
    .B(_13235_),
    .C(_13222_),
    .Y(_13236_));
 sky130_fd_sc_hd__a21oi_4 _35591_ (.A1(_12920_),
    .A2(_12919_),
    .B1(_12923_),
    .Y(_13237_));
 sky130_vsdinv _35592_ (.A(_13237_),
    .Y(_13238_));
 sky130_fd_sc_hd__a21o_2 _35593_ (.A1(_13233_),
    .A2(_13236_),
    .B1(_13238_),
    .X(_13239_));
 sky130_fd_sc_hd__a31oi_4 _35594_ (.A1(_13234_),
    .A2(_13235_),
    .A3(_13222_),
    .B1(_13237_),
    .Y(_13240_));
 sky130_fd_sc_hd__nand2_4 _35595_ (.A(_13240_),
    .B(_13233_),
    .Y(_13241_));
 sky130_fd_sc_hd__o21ai_2 _35596_ (.A1(_12554_),
    .A2(_12930_),
    .B1(_12925_),
    .Y(_13242_));
 sky130_fd_sc_hd__nand2_1 _35597_ (.A(_13242_),
    .B(_12929_),
    .Y(_13243_));
 sky130_fd_sc_hd__a21boi_4 _35598_ (.A1(_13239_),
    .A2(_13241_),
    .B1_N(_13243_),
    .Y(_13244_));
 sky130_fd_sc_hd__a21oi_2 _35599_ (.A1(_13234_),
    .A2(_13235_),
    .B1(_13222_),
    .Y(_13245_));
 sky130_fd_sc_hd__nand2_1 _35600_ (.A(_13236_),
    .B(_13238_),
    .Y(_13246_));
 sky130_fd_sc_hd__o2111a_2 _35601_ (.A1(_13245_),
    .A2(_13246_),
    .B1(_12929_),
    .C1(_13242_),
    .D1(_13239_),
    .X(_13247_));
 sky130_fd_sc_hd__buf_6 _35602_ (.A(_09817_),
    .X(_13248_));
 sky130_fd_sc_hd__a22oi_4 _35603_ (.A1(_19653_),
    .A2(_13248_),
    .B1(_19656_),
    .B2(_19840_),
    .Y(_13249_));
 sky130_fd_sc_hd__and4_2 _35604_ (.A(_19653_),
    .B(_06160_),
    .C(_10601_),
    .D(_19844_),
    .X(_13250_));
 sky130_fd_sc_hd__nand2_2 _35605_ (.A(net456),
    .B(_12639_),
    .Y(_13251_));
 sky130_fd_sc_hd__o21ai_4 _35606_ (.A1(_13249_),
    .A2(_13250_),
    .B1(_13251_),
    .Y(_13252_));
 sky130_fd_sc_hd__nand2_1 _35607_ (.A(_19653_),
    .B(_19844_),
    .Y(_13253_));
 sky130_fd_sc_hd__nand3b_4 _35608_ (.A_N(_13253_),
    .B(_19656_),
    .C(_11583_),
    .Y(_13254_));
 sky130_vsdinv _35609_ (.A(_13251_),
    .Y(_13255_));
 sky130_fd_sc_hd__a22o_1 _35610_ (.A1(_19653_),
    .A2(_10493_),
    .B1(_19656_),
    .B2(_11574_),
    .X(_13256_));
 sky130_fd_sc_hd__nand3_4 _35611_ (.A(_13254_),
    .B(_13255_),
    .C(_13256_),
    .Y(_13257_));
 sky130_fd_sc_hd__nand2_8 _35612_ (.A(_13252_),
    .B(_13257_),
    .Y(_13258_));
 sky130_vsdinv _35613_ (.A(_13258_),
    .Y(_13259_));
 sky130_fd_sc_hd__buf_6 _35614_ (.A(_10617_),
    .X(_13260_));
 sky130_fd_sc_hd__nand2_2 _35615_ (.A(_19644_),
    .B(_08773_),
    .Y(_13261_));
 sky130_fd_sc_hd__a21o_1 _35616_ (.A1(_19648_),
    .A2(_11224_),
    .B1(_13261_),
    .X(_13262_));
 sky130_fd_sc_hd__nand2_2 _35617_ (.A(_06416_),
    .B(_08787_),
    .Y(_13263_));
 sky130_fd_sc_hd__a21o_1 _35618_ (.A1(_19645_),
    .A2(_19855_),
    .B1(_13263_),
    .X(_13264_));
 sky130_fd_sc_hd__o211ai_4 _35619_ (.A1(net473),
    .A2(_13260_),
    .B1(_13262_),
    .C1(_13264_),
    .Y(_13265_));
 sky130_fd_sc_hd__nand3_2 _35620_ (.A(_08597_),
    .B(_09439_),
    .C(_10643_),
    .Y(_13266_));
 sky130_fd_sc_hd__nand2_1 _35621_ (.A(_13261_),
    .B(_13263_),
    .Y(_13267_));
 sky130_fd_sc_hd__o2111ai_4 _35622_ (.A1(_11537_),
    .A2(_13266_),
    .B1(net478),
    .C1(_19849_),
    .D1(_13267_),
    .Y(_13268_));
 sky130_fd_sc_hd__a21o_1 _35623_ (.A1(_12890_),
    .A2(_12892_),
    .B1(_12889_),
    .X(_13269_));
 sky130_fd_sc_hd__a21o_1 _35624_ (.A1(_13265_),
    .A2(_13268_),
    .B1(_13269_),
    .X(_13270_));
 sky130_fd_sc_hd__nand3_4 _35625_ (.A(_13269_),
    .B(_13265_),
    .C(_13268_),
    .Y(_13271_));
 sky130_fd_sc_hd__nand2_4 _35626_ (.A(_13270_),
    .B(_13271_),
    .Y(_13272_));
 sky130_fd_sc_hd__xor2_4 _35627_ (.A(_13259_),
    .B(_13272_),
    .X(_13273_));
 sky130_fd_sc_hd__o21ai_2 _35628_ (.A1(_13244_),
    .A2(_13247_),
    .B1(_13273_),
    .Y(_13274_));
 sky130_fd_sc_hd__xor2_4 _35629_ (.A(_13258_),
    .B(_13272_),
    .X(_13275_));
 sky130_fd_sc_hd__a22o_2 _35630_ (.A1(_12929_),
    .A2(_13242_),
    .B1(_13239_),
    .B2(_13241_),
    .X(_13276_));
 sky130_fd_sc_hd__nand3b_4 _35631_ (.A_N(_13243_),
    .B(_13239_),
    .C(_13241_),
    .Y(_13277_));
 sky130_fd_sc_hd__nand3_4 _35632_ (.A(_13275_),
    .B(_13276_),
    .C(_13277_),
    .Y(_13278_));
 sky130_fd_sc_hd__nand3b_4 _35633_ (.A_N(_13220_),
    .B(_13274_),
    .C(_13278_),
    .Y(_13279_));
 sky130_fd_sc_hd__o21ai_4 _35634_ (.A1(_13244_),
    .A2(_13247_),
    .B1(_13275_),
    .Y(_13280_));
 sky130_fd_sc_hd__nand3_4 _35635_ (.A(_13273_),
    .B(_13276_),
    .C(_13277_),
    .Y(_13281_));
 sky130_fd_sc_hd__nand3_4 _35636_ (.A(_13280_),
    .B(_13220_),
    .C(_13281_),
    .Y(_13282_));
 sky130_fd_sc_hd__nor2_4 _35637_ (.A(_12944_),
    .B(_12935_),
    .Y(_13283_));
 sky130_fd_sc_hd__nor2_8 _35638_ (.A(_12938_),
    .B(_13283_),
    .Y(_13284_));
 sky130_fd_sc_hd__a21oi_1 _35639_ (.A1(_13279_),
    .A2(_13282_),
    .B1(_13284_),
    .Y(_13285_));
 sky130_fd_sc_hd__nand3_4 _35640_ (.A(_13279_),
    .B(_13282_),
    .C(_13284_),
    .Y(_13286_));
 sky130_vsdinv _35641_ (.A(_13286_),
    .Y(_13287_));
 sky130_fd_sc_hd__o2bb2ai_2 _35642_ (.A1_N(_13211_),
    .A2_N(_13219_),
    .B1(_13285_),
    .B2(_13287_),
    .Y(_13288_));
 sky130_vsdinv _35643_ (.A(_13284_),
    .Y(_13289_));
 sky130_fd_sc_hd__a21oi_4 _35644_ (.A1(_13279_),
    .A2(_13282_),
    .B1(_13289_),
    .Y(_13290_));
 sky130_fd_sc_hd__and3_1 _35645_ (.A(_13279_),
    .B(_13289_),
    .C(_13282_),
    .X(_13291_));
 sky130_fd_sc_hd__o211ai_2 _35646_ (.A1(_13290_),
    .A2(_13291_),
    .B1(_13211_),
    .C1(_13219_),
    .Y(_13292_));
 sky130_fd_sc_hd__nand3_4 _35647_ (.A(_13092_),
    .B(_13288_),
    .C(_13292_),
    .Y(_13293_));
 sky130_fd_sc_hd__a21oi_1 _35648_ (.A1(_12870_),
    .A2(_12876_),
    .B1(_12874_),
    .Y(_13294_));
 sky130_fd_sc_hd__o21ai_2 _35649_ (.A1(_12966_),
    .A2(_13294_),
    .B1(_12877_),
    .Y(_13295_));
 sky130_fd_sc_hd__o2bb2ai_2 _35650_ (.A1_N(_13211_),
    .A2_N(_13219_),
    .B1(_13291_),
    .B2(_13290_),
    .Y(_13296_));
 sky130_fd_sc_hd__a21o_1 _35651_ (.A1(_13279_),
    .A2(_13282_),
    .B1(_13284_),
    .X(_13297_));
 sky130_fd_sc_hd__nand2_4 _35652_ (.A(_13297_),
    .B(_13286_),
    .Y(_13298_));
 sky130_fd_sc_hd__nand3_4 _35653_ (.A(_13298_),
    .B(_13211_),
    .C(_13219_),
    .Y(_13299_));
 sky130_fd_sc_hd__nand3_4 _35654_ (.A(_13295_),
    .B(_13296_),
    .C(_13299_),
    .Y(_13300_));
 sky130_fd_sc_hd__nand2_2 _35655_ (.A(_12904_),
    .B(_12905_),
    .Y(_13301_));
 sky130_fd_sc_hd__a21oi_4 _35656_ (.A1(_12909_),
    .A2(_13301_),
    .B1(_12906_),
    .Y(_13302_));
 sky130_fd_sc_hd__a22oi_4 _35657_ (.A1(_06493_),
    .A2(_11199_),
    .B1(_06505_),
    .B2(_11200_),
    .Y(_13303_));
 sky130_fd_sc_hd__nand3_4 _35658_ (.A(_05841_),
    .B(_19665_),
    .C(_19825_),
    .Y(_13304_));
 sky130_fd_sc_hd__nor2_2 _35659_ (.A(_10597_),
    .B(_13304_),
    .Y(_13305_));
 sky130_fd_sc_hd__nand2_4 _35660_ (.A(_18467_),
    .B(\pcpi_mul.rs2[6] ),
    .Y(_13306_));
 sky130_fd_sc_hd__clkinv_4 _35661_ (.A(_13306_),
    .Y(_13307_));
 sky130_fd_sc_hd__o21ai_2 _35662_ (.A1(_13303_),
    .A2(_13305_),
    .B1(_13307_),
    .Y(_13308_));
 sky130_fd_sc_hd__buf_6 _35663_ (.A(_10596_),
    .X(_13309_));
 sky130_fd_sc_hd__buf_4 _35664_ (.A(_13306_),
    .X(_13310_));
 sky130_fd_sc_hd__a22o_2 _35665_ (.A1(_05452_),
    .A2(_11199_),
    .B1(_05405_),
    .B2(_11597_),
    .X(_13311_));
 sky130_fd_sc_hd__o211ai_4 _35666_ (.A1(_13309_),
    .A2(_13304_),
    .B1(_13310_),
    .C1(_13311_),
    .Y(_13312_));
 sky130_fd_sc_hd__nand3_4 _35667_ (.A(_13302_),
    .B(_13308_),
    .C(_13312_),
    .Y(_13313_));
 sky130_fd_sc_hd__a31o_1 _35668_ (.A1(_13301_),
    .A2(net456),
    .A3(_19840_),
    .B1(_12906_),
    .X(_13314_));
 sky130_fd_sc_hd__o21ai_2 _35669_ (.A1(_13303_),
    .A2(_13305_),
    .B1(_13310_),
    .Y(_13315_));
 sky130_fd_sc_hd__o211ai_4 _35670_ (.A1(_13309_),
    .A2(_13304_),
    .B1(_13307_),
    .C1(_13311_),
    .Y(_13316_));
 sky130_fd_sc_hd__nand3_4 _35671_ (.A(_13314_),
    .B(_13315_),
    .C(_13316_),
    .Y(_13317_));
 sky130_fd_sc_hd__nor2_4 _35672_ (.A(_12977_),
    .B(_12970_),
    .Y(_13318_));
 sky130_fd_sc_hd__o2bb2ai_4 _35673_ (.A1_N(_13313_),
    .A2_N(_13317_),
    .B1(_12976_),
    .B2(_13318_),
    .Y(_13319_));
 sky130_fd_sc_hd__nor2_2 _35674_ (.A(_12976_),
    .B(_13318_),
    .Y(_13320_));
 sky130_fd_sc_hd__nand3_4 _35675_ (.A(_13317_),
    .B(_13313_),
    .C(_13320_),
    .Y(_13321_));
 sky130_vsdinv _35676_ (.A(_12893_),
    .Y(_13322_));
 sky130_fd_sc_hd__nand2_1 _35677_ (.A(_12888_),
    .B(_12895_),
    .Y(_13323_));
 sky130_fd_sc_hd__o2bb2ai_4 _35678_ (.A1_N(_12900_),
    .A2_N(_12911_),
    .B1(_13322_),
    .B2(_13323_),
    .Y(_13324_));
 sky130_fd_sc_hd__a21oi_4 _35679_ (.A1(_13319_),
    .A2(_13321_),
    .B1(_13324_),
    .Y(_13325_));
 sky130_fd_sc_hd__and3_1 _35680_ (.A(_13314_),
    .B(_13315_),
    .C(_13316_),
    .X(_13326_));
 sky130_fd_sc_hd__nand2_1 _35681_ (.A(_13313_),
    .B(_13320_),
    .Y(_13327_));
 sky130_fd_sc_hd__o211a_2 _35682_ (.A1(_13326_),
    .A2(_13327_),
    .B1(_13319_),
    .C1(_13324_),
    .X(_13328_));
 sky130_fd_sc_hd__nand2_1 _35683_ (.A(_12979_),
    .B(_12984_),
    .Y(_13329_));
 sky130_fd_sc_hd__nand2_4 _35684_ (.A(_13329_),
    .B(_12983_),
    .Y(_13330_));
 sky130_fd_sc_hd__o21ai_2 _35685_ (.A1(_13325_),
    .A2(_13328_),
    .B1(_13330_),
    .Y(_13331_));
 sky130_fd_sc_hd__a21boi_2 _35686_ (.A1(_12988_),
    .A2(_12996_),
    .B1_N(_12992_),
    .Y(_13332_));
 sky130_fd_sc_hd__a21o_1 _35687_ (.A1(_13319_),
    .A2(_13321_),
    .B1(_13324_),
    .X(_13333_));
 sky130_fd_sc_hd__nand3_2 _35688_ (.A(_13324_),
    .B(_13319_),
    .C(_13321_),
    .Y(_13334_));
 sky130_vsdinv _35689_ (.A(_13330_),
    .Y(_13335_));
 sky130_fd_sc_hd__nand3_2 _35690_ (.A(_13333_),
    .B(_13334_),
    .C(_13335_),
    .Y(_13336_));
 sky130_fd_sc_hd__nand3_4 _35691_ (.A(_13331_),
    .B(_13332_),
    .C(_13336_),
    .Y(_13337_));
 sky130_fd_sc_hd__o21ai_2 _35692_ (.A1(_13325_),
    .A2(_13328_),
    .B1(_13335_),
    .Y(_13338_));
 sky130_fd_sc_hd__nand2_1 _35693_ (.A(_12989_),
    .B(_12991_),
    .Y(_13339_));
 sky130_fd_sc_hd__a21oi_2 _35694_ (.A1(_12991_),
    .A2(_12990_),
    .B1(_12989_),
    .Y(_13340_));
 sky130_fd_sc_hd__o22ai_4 _35695_ (.A1(_12986_),
    .A2(_13339_),
    .B1(_12994_),
    .B2(_13340_),
    .Y(_13341_));
 sky130_fd_sc_hd__nand3_2 _35696_ (.A(_13333_),
    .B(_13334_),
    .C(_13330_),
    .Y(_13342_));
 sky130_fd_sc_hd__nand3_4 _35697_ (.A(_13338_),
    .B(_13341_),
    .C(_13342_),
    .Y(_13343_));
 sky130_fd_sc_hd__nand2_1 _35698_ (.A(_13337_),
    .B(_13343_),
    .Y(_13344_));
 sky130_fd_sc_hd__nand2_2 _35699_ (.A(_12279_),
    .B(_13005_),
    .Y(_13345_));
 sky130_fd_sc_hd__nand3_1 _35700_ (.A(_12281_),
    .B(_13004_),
    .C(_13009_),
    .Y(_13346_));
 sky130_fd_sc_hd__nand2_1 _35701_ (.A(_13345_),
    .B(_13346_),
    .Y(_13347_));
 sky130_fd_sc_hd__or2_2 _35702_ (.A(_12633_),
    .B(_13347_),
    .X(_13348_));
 sky130_fd_sc_hd__nand2_1 _35703_ (.A(_13347_),
    .B(_12633_),
    .Y(_13349_));
 sky130_fd_sc_hd__nand2_2 _35704_ (.A(_13348_),
    .B(_13349_),
    .Y(_13350_));
 sky130_fd_sc_hd__nand2_1 _35705_ (.A(_13344_),
    .B(_13350_),
    .Y(_13351_));
 sky130_vsdinv _35706_ (.A(_12949_),
    .Y(_13352_));
 sky130_fd_sc_hd__nand2_1 _35707_ (.A(_12947_),
    .B(_12950_),
    .Y(_13353_));
 sky130_fd_sc_hd__o2bb2ai_2 _35708_ (.A1_N(_12946_),
    .A2_N(_12952_),
    .B1(_13352_),
    .B2(_13353_),
    .Y(_13354_));
 sky130_vsdinv _35709_ (.A(_13350_),
    .Y(_13355_));
 sky130_fd_sc_hd__nand3_2 _35710_ (.A(_13355_),
    .B(_13337_),
    .C(_13343_),
    .Y(_13356_));
 sky130_fd_sc_hd__nand3_4 _35711_ (.A(_13351_),
    .B(_13354_),
    .C(_13356_),
    .Y(_13357_));
 sky130_fd_sc_hd__nand2_1 _35712_ (.A(_13344_),
    .B(_13355_),
    .Y(_13358_));
 sky130_fd_sc_hd__a21oi_4 _35713_ (.A1(_12946_),
    .A2(_12952_),
    .B1(_12963_),
    .Y(_13359_));
 sky130_fd_sc_hd__nand3_2 _35714_ (.A(_13337_),
    .B(_13343_),
    .C(_13350_),
    .Y(_13360_));
 sky130_fd_sc_hd__nand3_4 _35715_ (.A(_13358_),
    .B(_13359_),
    .C(_13360_),
    .Y(_13361_));
 sky130_fd_sc_hd__nand2_4 _35716_ (.A(_13027_),
    .B(_13000_),
    .Y(_13362_));
 sky130_fd_sc_hd__a21oi_4 _35717_ (.A1(_13357_),
    .A2(_13361_),
    .B1(_13362_),
    .Y(_13363_));
 sky130_fd_sc_hd__nand3_4 _35718_ (.A(_13357_),
    .B(_13361_),
    .C(_13362_),
    .Y(_13364_));
 sky130_vsdinv _35719_ (.A(_13364_),
    .Y(_13365_));
 sky130_fd_sc_hd__o2bb2ai_4 _35720_ (.A1_N(_13293_),
    .A2_N(_13300_),
    .B1(_13363_),
    .B2(_13365_),
    .Y(_13366_));
 sky130_fd_sc_hd__nor2_4 _35721_ (.A(_13363_),
    .B(_13365_),
    .Y(_13367_));
 sky130_fd_sc_hd__nand3_4 _35722_ (.A(_13367_),
    .B(_13300_),
    .C(_13293_),
    .Y(_13368_));
 sky130_fd_sc_hd__nand2_4 _35723_ (.A(_13046_),
    .B(_12958_),
    .Y(_13369_));
 sky130_fd_sc_hd__a21oi_4 _35724_ (.A1(_13366_),
    .A2(_13368_),
    .B1(_13369_),
    .Y(_13370_));
 sky130_fd_sc_hd__nand2_1 _35725_ (.A(_13296_),
    .B(_13299_),
    .Y(_13371_));
 sky130_fd_sc_hd__nand2_1 _35726_ (.A(_13357_),
    .B(_13361_),
    .Y(_13372_));
 sky130_fd_sc_hd__nor2_1 _35727_ (.A(_13021_),
    .B(_13022_),
    .Y(_13373_));
 sky130_fd_sc_hd__nand2_1 _35728_ (.A(_13372_),
    .B(_13373_),
    .Y(_13374_));
 sky130_fd_sc_hd__nand2_1 _35729_ (.A(_13374_),
    .B(_13364_),
    .Y(_13375_));
 sky130_fd_sc_hd__a21oi_1 _35730_ (.A1(_13371_),
    .A2(_13092_),
    .B1(_13375_),
    .Y(_13376_));
 sky130_fd_sc_hd__a2bb2oi_1 _35731_ (.A1_N(_13363_),
    .A2_N(_13365_),
    .B1(_13293_),
    .B2(_13300_),
    .Y(_13377_));
 sky130_fd_sc_hd__a221oi_2 _35732_ (.A1(_13046_),
    .A2(_12958_),
    .B1(_13376_),
    .B2(_13300_),
    .C1(_13377_),
    .Y(_13378_));
 sky130_fd_sc_hd__o22ai_4 _35733_ (.A1(_13089_),
    .A2(_13091_),
    .B1(_13370_),
    .B2(_13378_),
    .Y(_13379_));
 sky130_fd_sc_hd__a21o_1 _35734_ (.A1(_13366_),
    .A2(_13368_),
    .B1(_13369_),
    .X(_13380_));
 sky130_fd_sc_hd__nand3_4 _35735_ (.A(_13369_),
    .B(_13366_),
    .C(_13368_),
    .Y(_13381_));
 sky130_fd_sc_hd__xor2_4 _35736_ (.A(_13090_),
    .B(_13087_),
    .X(_13382_));
 sky130_fd_sc_hd__nand3_4 _35737_ (.A(_13380_),
    .B(_13381_),
    .C(_13382_),
    .Y(_13383_));
 sky130_fd_sc_hd__nand3_4 _35738_ (.A(_13084_),
    .B(_13379_),
    .C(_13383_),
    .Y(_13384_));
 sky130_fd_sc_hd__nor2_8 _35739_ (.A(_13090_),
    .B(_13088_),
    .Y(_13385_));
 sky130_fd_sc_hd__nor2_2 _35740_ (.A(_13086_),
    .B(_13087_),
    .Y(_13386_));
 sky130_fd_sc_hd__o22ai_4 _35741_ (.A1(_13385_),
    .A2(_13386_),
    .B1(_13370_),
    .B2(_13378_),
    .Y(_13387_));
 sky130_fd_sc_hd__o21ai_2 _35742_ (.A1(_13062_),
    .A2(_13043_),
    .B1(_13061_),
    .Y(_13388_));
 sky130_fd_sc_hd__nand3b_4 _35743_ (.A_N(_13382_),
    .B(_13380_),
    .C(_13381_),
    .Y(_13389_));
 sky130_fd_sc_hd__nand3_4 _35744_ (.A(_13387_),
    .B(_13388_),
    .C(_13389_),
    .Y(_13390_));
 sky130_fd_sc_hd__and3_2 _35745_ (.A(_13384_),
    .B(_13390_),
    .C(_13065_),
    .X(_13391_));
 sky130_vsdinv _35746_ (.A(_13065_),
    .Y(_13392_));
 sky130_fd_sc_hd__nand2_1 _35747_ (.A(_13384_),
    .B(_13390_),
    .Y(_13393_));
 sky130_fd_sc_hd__and3_1 _35748_ (.A(_13066_),
    .B(_13067_),
    .C(_13068_),
    .X(_13394_));
 sky130_fd_sc_hd__o2bb2ai_2 _35749_ (.A1_N(_13392_),
    .A2_N(_13393_),
    .B1(_13394_),
    .B2(_13077_),
    .Y(_13395_));
 sky130_fd_sc_hd__nor2_1 _35750_ (.A(_13391_),
    .B(_13395_),
    .Y(_13396_));
 sky130_vsdinv _35751_ (.A(_13396_),
    .Y(_13397_));
 sky130_fd_sc_hd__a21oi_2 _35752_ (.A1(_13384_),
    .A2(_13390_),
    .B1(_13065_),
    .Y(_13398_));
 sky130_fd_sc_hd__nor2_2 _35753_ (.A(_13394_),
    .B(_13077_),
    .Y(_13399_));
 sky130_fd_sc_hd__o21ai_4 _35754_ (.A1(_13398_),
    .A2(_13391_),
    .B1(_13399_),
    .Y(_13400_));
 sky130_fd_sc_hd__nand2_2 _35755_ (.A(_13397_),
    .B(_13400_),
    .Y(_13401_));
 sky130_fd_sc_hd__o2bb2ai_2 _35756_ (.A1_N(_12723_),
    .A2_N(_13079_),
    .B1(_13072_),
    .B2(_13074_),
    .Y(_13402_));
 sky130_fd_sc_hd__o2111ai_4 _35757_ (.A1(_13071_),
    .A2(_13402_),
    .B1(_12738_),
    .C1(_13076_),
    .D1(_12735_),
    .Y(_13403_));
 sky130_fd_sc_hd__or2_1 _35758_ (.A(_13403_),
    .B(_12748_),
    .X(_13404_));
 sky130_fd_sc_hd__nand2_1 _35759_ (.A(_12738_),
    .B(_13081_),
    .Y(_13405_));
 sky130_fd_sc_hd__nand2_2 _35760_ (.A(_13405_),
    .B(_13076_),
    .Y(_13406_));
 sky130_fd_sc_hd__nand2_2 _35761_ (.A(_13404_),
    .B(_13406_),
    .Y(_13407_));
 sky130_fd_sc_hd__xnor2_4 _35762_ (.A(_13401_),
    .B(_13407_),
    .Y(_02657_));
 sky130_fd_sc_hd__buf_4 _35763_ (.A(_19628_),
    .X(_13408_));
 sky130_fd_sc_hd__nor2_2 _35764_ (.A(_13186_),
    .B(_13187_),
    .Y(_13409_));
 sky130_fd_sc_hd__a31o_1 _35765_ (.A1(_13189_),
    .A2(_13408_),
    .A3(_19870_),
    .B1(_13409_),
    .X(_13410_));
 sky130_fd_sc_hd__nand3_4 _35766_ (.A(_19632_),
    .B(_19636_),
    .C(_08332_),
    .Y(_13411_));
 sky130_fd_sc_hd__nor2_8 _35767_ (.A(_10466_),
    .B(_13411_),
    .Y(_13412_));
 sky130_fd_sc_hd__buf_4 _35768_ (.A(_10453_),
    .X(_13413_));
 sky130_fd_sc_hd__a22o_2 _35769_ (.A1(_19633_),
    .A2(_10981_),
    .B1(_19637_),
    .B2(_13413_),
    .X(_13414_));
 sky130_fd_sc_hd__nand2_4 _35770_ (.A(_07435_),
    .B(_11232_),
    .Y(_13415_));
 sky130_vsdinv _35771_ (.A(_13415_),
    .Y(_13416_));
 sky130_fd_sc_hd__nand3b_2 _35772_ (.A_N(_13412_),
    .B(_13414_),
    .C(_13416_),
    .Y(_13417_));
 sky130_fd_sc_hd__a22oi_4 _35773_ (.A1(_10990_),
    .A2(_10981_),
    .B1(_10991_),
    .B2(_19859_),
    .Y(_13418_));
 sky130_fd_sc_hd__o21ai_2 _35774_ (.A1(_13418_),
    .A2(_13412_),
    .B1(_13415_),
    .Y(_13419_));
 sky130_fd_sc_hd__nand3_4 _35775_ (.A(_13410_),
    .B(_13417_),
    .C(_13419_),
    .Y(_13420_));
 sky130_fd_sc_hd__nand3b_2 _35776_ (.A_N(_13412_),
    .B(_13414_),
    .C(_13415_),
    .Y(_13421_));
 sky130_fd_sc_hd__a31oi_4 _35777_ (.A1(_13189_),
    .A2(_13408_),
    .A3(_19870_),
    .B1(_13409_),
    .Y(_13422_));
 sky130_fd_sc_hd__o21ai_2 _35778_ (.A1(_13418_),
    .A2(_13412_),
    .B1(_13416_),
    .Y(_13423_));
 sky130_fd_sc_hd__nand3_4 _35779_ (.A(_13421_),
    .B(_13422_),
    .C(_13423_),
    .Y(_13424_));
 sky130_fd_sc_hd__nor2_4 _35780_ (.A(_13231_),
    .B(_13225_),
    .Y(_13425_));
 sky130_fd_sc_hd__o2bb2ai_4 _35781_ (.A1_N(_13420_),
    .A2_N(_13424_),
    .B1(_13226_),
    .B2(_13425_),
    .Y(_13426_));
 sky130_fd_sc_hd__nor2_4 _35782_ (.A(_13226_),
    .B(_13425_),
    .Y(_13427_));
 sky130_fd_sc_hd__nand3_4 _35783_ (.A(_13420_),
    .B(_13424_),
    .C(_13427_),
    .Y(_13428_));
 sky130_fd_sc_hd__nand2_2 _35784_ (.A(_13246_),
    .B(_13233_),
    .Y(_13429_));
 sky130_fd_sc_hd__a21oi_2 _35785_ (.A1(_13426_),
    .A2(_13428_),
    .B1(_13429_),
    .Y(_13430_));
 sky130_fd_sc_hd__o211a_1 _35786_ (.A1(_13245_),
    .A2(_13240_),
    .B1(_13428_),
    .C1(_13426_),
    .X(_13431_));
 sky130_fd_sc_hd__a22oi_4 _35787_ (.A1(net445),
    .A2(_09823_),
    .B1(_06423_),
    .B2(_11909_),
    .Y(_13432_));
 sky130_fd_sc_hd__nand3_4 _35788_ (.A(_06606_),
    .B(_06907_),
    .C(_19851_),
    .Y(_13433_));
 sky130_fd_sc_hd__nor2_4 _35789_ (.A(_10617_),
    .B(_13433_),
    .Y(_13434_));
 sky130_fd_sc_hd__o22ai_4 _35790_ (.A1(net473),
    .A2(_10497_),
    .B1(_13432_),
    .B2(_13434_),
    .Y(_13435_));
 sky130_fd_sc_hd__a22o_1 _35791_ (.A1(_08597_),
    .A2(_19851_),
    .B1(_09439_),
    .B2(_11228_),
    .X(_13436_));
 sky130_fd_sc_hd__nor2_4 _35792_ (.A(_11721_),
    .B(_10496_),
    .Y(_13437_));
 sky130_fd_sc_hd__o211ai_4 _35793_ (.A1(_13260_),
    .A2(_13433_),
    .B1(_13436_),
    .C1(_13437_),
    .Y(_13438_));
 sky130_fd_sc_hd__o21ai_2 _35794_ (.A1(_13261_),
    .A2(_13263_),
    .B1(_13268_),
    .Y(_13439_));
 sky130_fd_sc_hd__a21oi_4 _35795_ (.A1(_13435_),
    .A2(_13438_),
    .B1(_13439_),
    .Y(_13440_));
 sky130_fd_sc_hd__nand2_1 _35796_ (.A(_13435_),
    .B(_13438_),
    .Y(_13441_));
 sky130_fd_sc_hd__o21a_1 _35797_ (.A1(_13261_),
    .A2(_13263_),
    .B1(_13268_),
    .X(_13442_));
 sky130_fd_sc_hd__nor2_2 _35798_ (.A(_13441_),
    .B(_13442_),
    .Y(_13443_));
 sky130_fd_sc_hd__a22oi_4 _35799_ (.A1(_06398_),
    .A2(_19839_),
    .B1(_06838_),
    .B2(_10598_),
    .Y(_13444_));
 sky130_fd_sc_hd__and4_2 _35800_ (.A(_06398_),
    .B(_06399_),
    .C(_10487_),
    .D(_09946_),
    .X(_13445_));
 sky130_fd_sc_hd__nor2_1 _35801_ (.A(_13444_),
    .B(_13445_),
    .Y(_13446_));
 sky130_fd_sc_hd__nand2_2 _35802_ (.A(_19659_),
    .B(_19829_),
    .Y(_13447_));
 sky130_fd_sc_hd__nand2_1 _35803_ (.A(_13446_),
    .B(_13447_),
    .Y(_13448_));
 sky130_vsdinv _35804_ (.A(_13447_),
    .Y(_13449_));
 sky130_fd_sc_hd__o21ai_1 _35805_ (.A1(_13444_),
    .A2(_13445_),
    .B1(_13449_),
    .Y(_13450_));
 sky130_fd_sc_hd__nand2_2 _35806_ (.A(_13448_),
    .B(_13450_),
    .Y(_13451_));
 sky130_fd_sc_hd__o21ai_1 _35807_ (.A1(_13440_),
    .A2(_13443_),
    .B1(_13451_),
    .Y(_13452_));
 sky130_vsdinv _35808_ (.A(_13435_),
    .Y(_13453_));
 sky130_fd_sc_hd__nand2_2 _35809_ (.A(_13439_),
    .B(_13438_),
    .Y(_13454_));
 sky130_fd_sc_hd__nand2_2 _35810_ (.A(_13442_),
    .B(_13441_),
    .Y(_13455_));
 sky130_fd_sc_hd__nand2_1 _35811_ (.A(_13446_),
    .B(_13449_),
    .Y(_13456_));
 sky130_fd_sc_hd__o21ai_1 _35812_ (.A1(_13444_),
    .A2(_13445_),
    .B1(_13447_),
    .Y(_13457_));
 sky130_fd_sc_hd__nand2_2 _35813_ (.A(_13456_),
    .B(_13457_),
    .Y(_13458_));
 sky130_fd_sc_hd__o211ai_2 _35814_ (.A1(_13453_),
    .A2(_13454_),
    .B1(_13455_),
    .C1(_13458_),
    .Y(_13459_));
 sky130_fd_sc_hd__nand2_2 _35815_ (.A(_13452_),
    .B(_13459_),
    .Y(_13460_));
 sky130_fd_sc_hd__o21bai_4 _35816_ (.A1(_13430_),
    .A2(_13431_),
    .B1_N(_13460_),
    .Y(_13461_));
 sky130_fd_sc_hd__a21o_1 _35817_ (.A1(_13426_),
    .A2(_13428_),
    .B1(_13429_),
    .X(_13462_));
 sky130_fd_sc_hd__nand3_4 _35818_ (.A(_13429_),
    .B(_13426_),
    .C(_13428_),
    .Y(_13463_));
 sky130_fd_sc_hd__nand3_4 _35819_ (.A(_13462_),
    .B(_13463_),
    .C(_13460_),
    .Y(_13464_));
 sky130_fd_sc_hd__o21ai_4 _35820_ (.A1(_13204_),
    .A2(_13203_),
    .B1(_13201_),
    .Y(_13465_));
 sky130_fd_sc_hd__a21o_1 _35821_ (.A1(_13461_),
    .A2(_13464_),
    .B1(_13465_),
    .X(_13466_));
 sky130_fd_sc_hd__nand3_4 _35822_ (.A(_13461_),
    .B(_13465_),
    .C(_13464_),
    .Y(_13467_));
 sky130_fd_sc_hd__a21oi_4 _35823_ (.A1(_13275_),
    .A2(_13276_),
    .B1(_13247_),
    .Y(_13468_));
 sky130_fd_sc_hd__a21boi_4 _35824_ (.A1(_13466_),
    .A2(_13467_),
    .B1_N(_13468_),
    .Y(_13469_));
 sky130_fd_sc_hd__a21oi_4 _35825_ (.A1(_13461_),
    .A2(_13464_),
    .B1(_13465_),
    .Y(_13470_));
 sky130_fd_sc_hd__nor2_2 _35826_ (.A(_13468_),
    .B(_13470_),
    .Y(_13471_));
 sky130_fd_sc_hd__nand2_1 _35827_ (.A(_13471_),
    .B(_13467_),
    .Y(_13472_));
 sky130_vsdinv _35828_ (.A(_13472_),
    .Y(_13473_));
 sky130_fd_sc_hd__nand3_4 _35829_ (.A(_08152_),
    .B(_19611_),
    .C(net497),
    .Y(_13474_));
 sky130_fd_sc_hd__nor2_8 _35830_ (.A(_07560_),
    .B(_13474_),
    .Y(_13475_));
 sky130_fd_sc_hd__nand2_4 _35831_ (.A(_19616_),
    .B(_07067_),
    .Y(_13476_));
 sky130_vsdinv _35832_ (.A(_13476_),
    .Y(_13477_));
 sky130_fd_sc_hd__a22o_2 _35833_ (.A1(_08153_),
    .A2(_19881_),
    .B1(_08155_),
    .B2(_08734_),
    .X(_13478_));
 sky130_fd_sc_hd__nand3b_2 _35834_ (.A_N(_13475_),
    .B(_13477_),
    .C(_13478_),
    .Y(_13479_));
 sky130_fd_sc_hd__a21o_1 _35835_ (.A1(_13177_),
    .A2(_13176_),
    .B1(_13172_),
    .X(_13480_));
 sky130_fd_sc_hd__a22oi_4 _35836_ (.A1(_08153_),
    .A2(_19881_),
    .B1(_08155_),
    .B2(_19878_),
    .Y(_13481_));
 sky130_fd_sc_hd__o21ai_2 _35837_ (.A1(_13481_),
    .A2(_13475_),
    .B1(_13476_),
    .Y(_13482_));
 sky130_fd_sc_hd__nand3_4 _35838_ (.A(_13479_),
    .B(_13480_),
    .C(_13482_),
    .Y(_13483_));
 sky130_fd_sc_hd__o21ai_2 _35839_ (.A1(_13481_),
    .A2(_13475_),
    .B1(_13477_),
    .Y(_13484_));
 sky130_fd_sc_hd__a21oi_4 _35840_ (.A1(_13177_),
    .A2(_13176_),
    .B1(_13172_),
    .Y(_13485_));
 sky130_fd_sc_hd__o211ai_4 _35841_ (.A1(_08447_),
    .A2(_13474_),
    .B1(_13476_),
    .C1(_13478_),
    .Y(_13486_));
 sky130_fd_sc_hd__nand3_4 _35842_ (.A(_13484_),
    .B(_13485_),
    .C(_13486_),
    .Y(_13487_));
 sky130_fd_sc_hd__nand2_1 _35843_ (.A(_13483_),
    .B(_13487_),
    .Y(_13488_));
 sky130_fd_sc_hd__nand2_4 _35844_ (.A(_07486_),
    .B(_07702_),
    .Y(_13489_));
 sky130_fd_sc_hd__nand2_4 _35845_ (.A(_08174_),
    .B(_08485_),
    .Y(_13490_));
 sky130_fd_sc_hd__nor2_2 _35846_ (.A(_13489_),
    .B(_13490_),
    .Y(_13491_));
 sky130_fd_sc_hd__and2_1 _35847_ (.A(_13489_),
    .B(_13490_),
    .X(_13492_));
 sky130_fd_sc_hd__nand2_1 _35848_ (.A(_19628_),
    .B(_10738_),
    .Y(_13493_));
 sky130_fd_sc_hd__o21bai_4 _35849_ (.A1(_13491_),
    .A2(_13492_),
    .B1_N(_13493_),
    .Y(_13494_));
 sky130_fd_sc_hd__a211o_2 _35850_ (.A1(_11003_),
    .A2(_19867_),
    .B1(_13491_),
    .C1(_13492_),
    .X(_13495_));
 sky130_fd_sc_hd__nand3_4 _35851_ (.A(_13488_),
    .B(_13494_),
    .C(_13495_),
    .Y(_13496_));
 sky130_fd_sc_hd__nand2_2 _35852_ (.A(_13495_),
    .B(_13494_),
    .Y(_13497_));
 sky130_fd_sc_hd__nand3_4 _35853_ (.A(_13497_),
    .B(_13487_),
    .C(_13483_),
    .Y(_13498_));
 sky130_fd_sc_hd__nand2_1 _35854_ (.A(_13496_),
    .B(_13498_),
    .Y(_13499_));
 sky130_fd_sc_hd__nand2_1 _35855_ (.A(_13153_),
    .B(_13155_),
    .Y(_13500_));
 sky130_fd_sc_hd__and2_1 _35856_ (.A(_13500_),
    .B(_13150_),
    .X(_13501_));
 sky130_fd_sc_hd__nand2_2 _35857_ (.A(_13499_),
    .B(_13501_),
    .Y(_13502_));
 sky130_fd_sc_hd__nand2_2 _35858_ (.A(_13500_),
    .B(_13150_),
    .Y(_13503_));
 sky130_fd_sc_hd__nand3_2 _35859_ (.A(_13503_),
    .B(_13496_),
    .C(_13498_),
    .Y(_13504_));
 sky130_fd_sc_hd__nand2_1 _35860_ (.A(_13502_),
    .B(_13504_),
    .Y(_13505_));
 sky130_fd_sc_hd__nand2_1 _35861_ (.A(_13193_),
    .B(_13180_),
    .Y(_13506_));
 sky130_fd_sc_hd__nand2_1 _35862_ (.A(_13506_),
    .B(_13184_),
    .Y(_13507_));
 sky130_fd_sc_hd__clkbuf_2 _35863_ (.A(_13507_),
    .X(_13508_));
 sky130_fd_sc_hd__and2_1 _35864_ (.A(_13505_),
    .B(_13508_),
    .X(_13509_));
 sky130_fd_sc_hd__a21oi_2 _35865_ (.A1(_13499_),
    .A2(_13501_),
    .B1(_13507_),
    .Y(_13510_));
 sky130_fd_sc_hd__clkbuf_2 _35866_ (.A(_13504_),
    .X(_13511_));
 sky130_fd_sc_hd__nand2_2 _35867_ (.A(_13510_),
    .B(_13511_),
    .Y(_13512_));
 sky130_vsdinv _35868_ (.A(_13512_),
    .Y(_13513_));
 sky130_fd_sc_hd__buf_4 _35869_ (.A(_10256_),
    .X(_13514_));
 sky130_fd_sc_hd__nand3_1 _35870_ (.A(_13514_),
    .B(_08947_),
    .C(_06284_),
    .Y(_13515_));
 sky130_fd_sc_hd__nand2_2 _35871_ (.A(_09722_),
    .B(_07072_),
    .Y(_13516_));
 sky130_fd_sc_hd__nand2_2 _35872_ (.A(_10257_),
    .B(_07642_),
    .Y(_13517_));
 sky130_fd_sc_hd__nand2_2 _35873_ (.A(_13516_),
    .B(_13517_),
    .Y(_13518_));
 sky130_fd_sc_hd__nand2_2 _35874_ (.A(_11801_),
    .B(_06634_),
    .Y(_13519_));
 sky130_vsdinv _35875_ (.A(_13519_),
    .Y(_13520_));
 sky130_fd_sc_hd__o211a_1 _35876_ (.A1(_06810_),
    .A2(_13515_),
    .B1(_13518_),
    .C1(_13520_),
    .X(_13521_));
 sky130_fd_sc_hd__o21a_1 _35877_ (.A1(_13119_),
    .A2(_13117_),
    .B1(_13129_),
    .X(_13522_));
 sky130_fd_sc_hd__nor2_4 _35878_ (.A(_13516_),
    .B(_13517_),
    .Y(_13523_));
 sky130_fd_sc_hd__and2_1 _35879_ (.A(_13516_),
    .B(_13517_),
    .X(_13524_));
 sky130_fd_sc_hd__o21ai_2 _35880_ (.A1(_13523_),
    .A2(_13524_),
    .B1(_13519_),
    .Y(_13525_));
 sky130_fd_sc_hd__nand3b_4 _35881_ (.A_N(_13521_),
    .B(_13522_),
    .C(_13525_),
    .Y(_13526_));
 sky130_fd_sc_hd__o21ai_2 _35882_ (.A1(_13523_),
    .A2(_13524_),
    .B1(_13520_),
    .Y(_13527_));
 sky130_fd_sc_hd__o21ai_2 _35883_ (.A1(_13119_),
    .A2(_13117_),
    .B1(_13129_),
    .Y(_13528_));
 sky130_fd_sc_hd__nand3b_2 _35884_ (.A_N(_13523_),
    .B(_13518_),
    .C(_13519_),
    .Y(_13529_));
 sky130_fd_sc_hd__nand3_4 _35885_ (.A(_13527_),
    .B(_13528_),
    .C(_13529_),
    .Y(_13530_));
 sky130_fd_sc_hd__a21oi_1 _35886_ (.A1(_13148_),
    .A2(_13147_),
    .B1(_13143_),
    .Y(_13531_));
 sky130_vsdinv _35887_ (.A(_13531_),
    .Y(_13532_));
 sky130_fd_sc_hd__a21oi_4 _35888_ (.A1(_13526_),
    .A2(_13530_),
    .B1(_13532_),
    .Y(_13533_));
 sky130_fd_sc_hd__nand3_4 _35889_ (.A(_13526_),
    .B(_13530_),
    .C(_13532_),
    .Y(_13534_));
 sky130_vsdinv _35890_ (.A(_13534_),
    .Y(_13535_));
 sky130_fd_sc_hd__a22oi_4 _35891_ (.A1(_19583_),
    .A2(_05811_),
    .B1(_10282_),
    .B2(_06119_),
    .Y(_13536_));
 sky130_fd_sc_hd__buf_2 _35892_ (.A(_13536_),
    .X(_13537_));
 sky130_fd_sc_hd__nand2_1 _35893_ (.A(_10281_),
    .B(_05804_),
    .Y(_13538_));
 sky130_fd_sc_hd__nand3b_4 _35894_ (.A_N(_13538_),
    .B(_19588_),
    .C(_10365_),
    .Y(_13539_));
 sky130_fd_sc_hd__nand2_4 _35895_ (.A(_10251_),
    .B(_06116_),
    .Y(_13540_));
 sky130_vsdinv _35896_ (.A(_13540_),
    .Y(_13541_));
 sky130_fd_sc_hd__nand2_1 _35897_ (.A(_13539_),
    .B(_13541_),
    .Y(_13542_));
 sky130_fd_sc_hd__nor2_2 _35898_ (.A(_13537_),
    .B(_13542_),
    .Y(_13543_));
 sky130_fd_sc_hd__and4_4 _35899_ (.A(_19583_),
    .B(_19588_),
    .C(_10365_),
    .D(_05799_),
    .X(_13544_));
 sky130_fd_sc_hd__o21ai_1 _35900_ (.A1(_13536_),
    .A2(_13544_),
    .B1(_13540_),
    .Y(_13545_));
 sky130_vsdinv _35901_ (.A(_13545_),
    .Y(_13546_));
 sky130_fd_sc_hd__o21ai_2 _35902_ (.A1(_13098_),
    .A2(_13105_),
    .B1(_13101_),
    .Y(_13547_));
 sky130_fd_sc_hd__nand3_4 _35903_ (.A(_12402_),
    .B(_12401_),
    .C(_06106_),
    .Y(_13548_));
 sky130_fd_sc_hd__nor2_4 _35904_ (.A(_19911_),
    .B(_13548_),
    .Y(_13549_));
 sky130_fd_sc_hd__a22oi_4 _35905_ (.A1(_12779_),
    .A2(_05808_),
    .B1(_06215_),
    .B2(_12781_),
    .Y(_13550_));
 sky130_fd_sc_hd__nand2_4 _35906_ (.A(net498),
    .B(_06827_),
    .Y(_13551_));
 sky130_fd_sc_hd__o21ai_4 _35907_ (.A1(_13549_),
    .A2(_13550_),
    .B1(_13551_),
    .Y(_13552_));
 sky130_fd_sc_hd__nand2_2 _35908_ (.A(_19576_),
    .B(_19907_),
    .Y(_13553_));
 sky130_fd_sc_hd__nand3b_4 _35909_ (.A_N(_13553_),
    .B(_13107_),
    .C(_06215_),
    .Y(_13554_));
 sky130_fd_sc_hd__o21ai_4 _35910_ (.A1(_19911_),
    .A2(_13099_),
    .B1(_13553_),
    .Y(_13555_));
 sky130_vsdinv _35911_ (.A(_13551_),
    .Y(_13556_));
 sky130_fd_sc_hd__nand3_4 _35912_ (.A(_13554_),
    .B(_13555_),
    .C(_13556_),
    .Y(_13557_));
 sky130_fd_sc_hd__a22oi_4 _35913_ (.A1(_13106_),
    .A2(_13547_),
    .B1(_13552_),
    .B2(_13557_),
    .Y(_13558_));
 sky130_fd_sc_hd__a21oi_4 _35914_ (.A1(_13105_),
    .A2(_13098_),
    .B1(_13101_),
    .Y(_13559_));
 sky130_fd_sc_hd__o211a_4 _35915_ (.A1(_13100_),
    .A2(_13559_),
    .B1(_13557_),
    .C1(_13552_),
    .X(_13560_));
 sky130_fd_sc_hd__o22ai_4 _35916_ (.A1(_13543_),
    .A2(_13546_),
    .B1(_13558_),
    .B2(_13560_),
    .Y(_13561_));
 sky130_fd_sc_hd__o21a_1 _35917_ (.A1(_13098_),
    .A2(_13105_),
    .B1(_13101_),
    .X(_13562_));
 sky130_fd_sc_hd__o21bai_1 _35918_ (.A1(_19911_),
    .A2(_13548_),
    .B1_N(_13551_),
    .Y(_13563_));
 sky130_fd_sc_hd__nor2_2 _35919_ (.A(_13550_),
    .B(_13563_),
    .Y(_13564_));
 sky130_fd_sc_hd__a21oi_2 _35920_ (.A1(_13554_),
    .A2(_13555_),
    .B1(_13556_),
    .Y(_13565_));
 sky130_fd_sc_hd__o22ai_4 _35921_ (.A1(_13097_),
    .A2(_13562_),
    .B1(_13564_),
    .B2(_13565_),
    .Y(_13566_));
 sky130_fd_sc_hd__o21a_2 _35922_ (.A1(_13537_),
    .A2(_13542_),
    .B1(_13545_),
    .X(_13567_));
 sky130_fd_sc_hd__o211ai_4 _35923_ (.A1(_13100_),
    .A2(_13559_),
    .B1(_13557_),
    .C1(_13552_),
    .Y(_13568_));
 sky130_fd_sc_hd__nand3_4 _35924_ (.A(_13566_),
    .B(_13567_),
    .C(_13568_),
    .Y(_13569_));
 sky130_vsdinv _35925_ (.A(_13113_),
    .Y(_13570_));
 sky130_fd_sc_hd__nand2_1 _35926_ (.A(_13111_),
    .B(_13112_),
    .Y(_13571_));
 sky130_fd_sc_hd__o2bb2ai_4 _35927_ (.A1_N(_13110_),
    .A2_N(_13137_),
    .B1(_13570_),
    .B2(_13571_),
    .Y(_13572_));
 sky130_fd_sc_hd__a21oi_4 _35928_ (.A1(_13561_),
    .A2(_13569_),
    .B1(_13572_),
    .Y(_13573_));
 sky130_fd_sc_hd__nand2_1 _35929_ (.A(_13566_),
    .B(_13567_),
    .Y(_13574_));
 sky130_fd_sc_hd__o211a_4 _35930_ (.A1(_13560_),
    .A2(_13574_),
    .B1(_13572_),
    .C1(_13561_),
    .X(_13575_));
 sky130_fd_sc_hd__o22ai_4 _35931_ (.A1(_13533_),
    .A2(_13535_),
    .B1(_13573_),
    .B2(_13575_),
    .Y(_13576_));
 sky130_fd_sc_hd__nor2_4 _35932_ (.A(_13533_),
    .B(_13535_),
    .Y(_13577_));
 sky130_fd_sc_hd__a21oi_2 _35933_ (.A1(_13566_),
    .A2(_13568_),
    .B1(_13567_),
    .Y(_13578_));
 sky130_fd_sc_hd__o21a_1 _35934_ (.A1(_13537_),
    .A2(_13544_),
    .B1(_13541_),
    .X(_13579_));
 sky130_fd_sc_hd__nor3_2 _35935_ (.A(_13541_),
    .B(_13537_),
    .C(_13544_),
    .Y(_13580_));
 sky130_fd_sc_hd__o211a_1 _35936_ (.A1(_13579_),
    .A2(_13580_),
    .B1(_13568_),
    .C1(_13566_),
    .X(_13581_));
 sky130_fd_sc_hd__o21bai_4 _35937_ (.A1(_13578_),
    .A2(_13581_),
    .B1_N(_13572_),
    .Y(_13582_));
 sky130_fd_sc_hd__nand3_4 _35938_ (.A(_13561_),
    .B(_13572_),
    .C(_13569_),
    .Y(_13583_));
 sky130_fd_sc_hd__nand3_4 _35939_ (.A(_13577_),
    .B(_13582_),
    .C(_13583_),
    .Y(_13584_));
 sky130_fd_sc_hd__nand2_1 _35940_ (.A(_13160_),
    .B(_13133_),
    .Y(_13585_));
 sky130_fd_sc_hd__nand2_4 _35941_ (.A(_13585_),
    .B(_13139_),
    .Y(_13586_));
 sky130_fd_sc_hd__a21oi_4 _35942_ (.A1(_13576_),
    .A2(_13584_),
    .B1(_13586_),
    .Y(_13587_));
 sky130_fd_sc_hd__and3_2 _35943_ (.A(_13576_),
    .B(_13586_),
    .C(_13584_),
    .X(_13588_));
 sky130_fd_sc_hd__o22ai_4 _35944_ (.A1(_13509_),
    .A2(_13513_),
    .B1(_13587_),
    .B2(_13588_),
    .Y(_13589_));
 sky130_fd_sc_hd__nand2_2 _35945_ (.A(_13505_),
    .B(_13508_),
    .Y(_13590_));
 sky130_fd_sc_hd__nand2_2 _35946_ (.A(_13590_),
    .B(_13512_),
    .Y(_13591_));
 sky130_fd_sc_hd__a21o_1 _35947_ (.A1(_13526_),
    .A2(_13530_),
    .B1(_13532_),
    .X(_13592_));
 sky130_fd_sc_hd__a22oi_4 _35948_ (.A1(_13592_),
    .A2(_13534_),
    .B1(_13582_),
    .B2(_13583_),
    .Y(_13593_));
 sky130_fd_sc_hd__nand2_2 _35949_ (.A(_13592_),
    .B(_13534_),
    .Y(_13594_));
 sky130_fd_sc_hd__nor3_4 _35950_ (.A(_13594_),
    .B(_13573_),
    .C(_13575_),
    .Y(_13595_));
 sky130_fd_sc_hd__o21bai_4 _35951_ (.A1(_13593_),
    .A2(_13595_),
    .B1_N(_13586_),
    .Y(_13596_));
 sky130_fd_sc_hd__nand3_4 _35952_ (.A(_13576_),
    .B(_13586_),
    .C(_13584_),
    .Y(_13597_));
 sky130_fd_sc_hd__nand3b_4 _35953_ (.A_N(_13591_),
    .B(_13596_),
    .C(_13597_),
    .Y(_13598_));
 sky130_fd_sc_hd__a21oi_4 _35954_ (.A1(_13158_),
    .A2(_13161_),
    .B1(_13096_),
    .Y(_13599_));
 sky130_fd_sc_hd__o21ai_4 _35955_ (.A1(_13599_),
    .A2(_13217_),
    .B1(_13162_),
    .Y(_13600_));
 sky130_fd_sc_hd__a21oi_4 _35956_ (.A1(_13589_),
    .A2(_13598_),
    .B1(_13600_),
    .Y(_13601_));
 sky130_vsdinv _35957_ (.A(_13162_),
    .Y(_13602_));
 sky130_fd_sc_hd__nor2_1 _35958_ (.A(_13599_),
    .B(_13217_),
    .Y(_13603_));
 sky130_fd_sc_hd__o211a_2 _35959_ (.A1(_13602_),
    .A2(_13603_),
    .B1(_13598_),
    .C1(_13589_),
    .X(_13604_));
 sky130_fd_sc_hd__o22ai_4 _35960_ (.A1(_13469_),
    .A2(_13473_),
    .B1(_13601_),
    .B2(_13604_),
    .Y(_13605_));
 sky130_fd_sc_hd__and3_1 _35961_ (.A(_13094_),
    .B(_13207_),
    .C(_13210_),
    .X(_13606_));
 sky130_fd_sc_hd__a21o_1 _35962_ (.A1(_13298_),
    .A2(_13219_),
    .B1(_13606_),
    .X(_13607_));
 sky130_fd_sc_hd__a22oi_4 _35963_ (.A1(_13590_),
    .A2(_13512_),
    .B1(_13596_),
    .B2(_13597_),
    .Y(_13608_));
 sky130_fd_sc_hd__nor3_4 _35964_ (.A(_13591_),
    .B(_13587_),
    .C(_13588_),
    .Y(_13609_));
 sky130_fd_sc_hd__o21bai_4 _35965_ (.A1(_13608_),
    .A2(_13609_),
    .B1_N(_13600_),
    .Y(_13610_));
 sky130_fd_sc_hd__nand3_4 _35966_ (.A(_13589_),
    .B(_13598_),
    .C(_13600_),
    .Y(_13611_));
 sky130_fd_sc_hd__a21oi_4 _35967_ (.A1(_13467_),
    .A2(_13471_),
    .B1(_13469_),
    .Y(_13612_));
 sky130_fd_sc_hd__nand3_4 _35968_ (.A(_13610_),
    .B(_13611_),
    .C(_13612_),
    .Y(_13613_));
 sky130_fd_sc_hd__nand3_4 _35969_ (.A(_13605_),
    .B(_13607_),
    .C(_13613_),
    .Y(_13614_));
 sky130_fd_sc_hd__o21ai_2 _35970_ (.A1(_13601_),
    .A2(_13604_),
    .B1(_13612_),
    .Y(_13615_));
 sky130_fd_sc_hd__a21oi_4 _35971_ (.A1(_13298_),
    .A2(_13219_),
    .B1(_13606_),
    .Y(_13616_));
 sky130_fd_sc_hd__nand2_1 _35972_ (.A(_13466_),
    .B(_13467_),
    .Y(_13617_));
 sky130_fd_sc_hd__nand2_1 _35973_ (.A(_13617_),
    .B(_13468_),
    .Y(_13618_));
 sky130_fd_sc_hd__nand2_2 _35974_ (.A(_13618_),
    .B(_13472_),
    .Y(_13619_));
 sky130_fd_sc_hd__nand3_4 _35975_ (.A(_13610_),
    .B(_13611_),
    .C(_13619_),
    .Y(_13620_));
 sky130_fd_sc_hd__nand3_4 _35976_ (.A(_13615_),
    .B(_13616_),
    .C(_13620_),
    .Y(_13621_));
 sky130_fd_sc_hd__a21oi_4 _35977_ (.A1(_13333_),
    .A2(_13330_),
    .B1(_13328_),
    .Y(_13622_));
 sky130_fd_sc_hd__a22oi_4 _35978_ (.A1(_11596_),
    .A2(_19666_),
    .B1(_19663_),
    .B2(_11200_),
    .Y(_13623_));
 sky130_fd_sc_hd__and4_1 _35979_ (.A(_11596_),
    .B(_06493_),
    .C(_06505_),
    .D(_11200_),
    .X(_13624_));
 sky130_fd_sc_hd__o21ai_2 _35980_ (.A1(_13623_),
    .A2(_13624_),
    .B1(_13307_),
    .Y(_13625_));
 sky130_fd_sc_hd__a21oi_2 _35981_ (.A1(_13256_),
    .A2(_13255_),
    .B1(_13250_),
    .Y(_13626_));
 sky130_fd_sc_hd__nand2_1 _35982_ (.A(_12614_),
    .B(_05843_),
    .Y(_13627_));
 sky130_fd_sc_hd__nand3b_4 _35983_ (.A_N(_13627_),
    .B(_19663_),
    .C(_19826_),
    .Y(_13628_));
 sky130_fd_sc_hd__a22o_1 _35984_ (.A1(_11594_),
    .A2(_19666_),
    .B1(_19663_),
    .B2(_19826_),
    .X(_13629_));
 sky130_fd_sc_hd__nand3_2 _35985_ (.A(_13628_),
    .B(_13310_),
    .C(_13629_),
    .Y(_13630_));
 sky130_fd_sc_hd__nand3_4 _35986_ (.A(_13625_),
    .B(_13626_),
    .C(_13630_),
    .Y(_13631_));
 sky130_fd_sc_hd__o21ai_2 _35987_ (.A1(_13623_),
    .A2(_13624_),
    .B1(_13310_),
    .Y(_13632_));
 sky130_fd_sc_hd__nand3_2 _35988_ (.A(_13628_),
    .B(_13307_),
    .C(_13629_),
    .Y(_13633_));
 sky130_fd_sc_hd__o21ai_2 _35989_ (.A1(_13251_),
    .A2(_13249_),
    .B1(_13254_),
    .Y(_13634_));
 sky130_fd_sc_hd__nand3_4 _35990_ (.A(_13632_),
    .B(_13633_),
    .C(_13634_),
    .Y(_13635_));
 sky130_fd_sc_hd__a21o_2 _35991_ (.A1(_13311_),
    .A2(_13307_),
    .B1(_13305_),
    .X(_13636_));
 sky130_fd_sc_hd__a21o_1 _35992_ (.A1(_13631_),
    .A2(_13635_),
    .B1(_13636_),
    .X(_13637_));
 sky130_fd_sc_hd__nand3_4 _35993_ (.A(_13631_),
    .B(_13635_),
    .C(_13636_),
    .Y(_13638_));
 sky130_fd_sc_hd__a21oi_2 _35994_ (.A1(_13265_),
    .A2(_13268_),
    .B1(_13269_),
    .Y(_13639_));
 sky130_fd_sc_hd__o21ai_4 _35995_ (.A1(_13258_),
    .A2(_13639_),
    .B1(_13271_),
    .Y(_13640_));
 sky130_fd_sc_hd__a21o_1 _35996_ (.A1(_13637_),
    .A2(_13638_),
    .B1(_13640_),
    .X(_13641_));
 sky130_fd_sc_hd__nand3_4 _35997_ (.A(_13640_),
    .B(_13637_),
    .C(_13638_),
    .Y(_13642_));
 sky130_fd_sc_hd__and2_2 _35998_ (.A(_13327_),
    .B(_13317_),
    .X(_13643_));
 sky130_fd_sc_hd__a21bo_1 _35999_ (.A1(_13641_),
    .A2(_13642_),
    .B1_N(_13643_),
    .X(_13644_));
 sky130_fd_sc_hd__nand3b_2 _36000_ (.A_N(_13643_),
    .B(_13641_),
    .C(_13642_),
    .Y(_13645_));
 sky130_fd_sc_hd__nand3b_4 _36001_ (.A_N(_13622_),
    .B(_13644_),
    .C(_13645_),
    .Y(_13646_));
 sky130_fd_sc_hd__a21o_1 _36002_ (.A1(_13641_),
    .A2(_13642_),
    .B1(_13643_),
    .X(_13647_));
 sky130_fd_sc_hd__nand3_2 _36003_ (.A(_13641_),
    .B(_13643_),
    .C(_13642_),
    .Y(_13648_));
 sky130_fd_sc_hd__nand3_4 _36004_ (.A(_13647_),
    .B(_13622_),
    .C(_13648_),
    .Y(_13649_));
 sky130_fd_sc_hd__a2111o_4 _36005_ (.A1(_12276_),
    .A2(_12277_),
    .B1(_12617_),
    .C1(_06447_),
    .D1(_11186_),
    .X(_13650_));
 sky130_fd_sc_hd__a21oi_4 _36006_ (.A1(_13650_),
    .A2(_13345_),
    .B1(_12635_),
    .Y(_13651_));
 sky130_fd_sc_hd__and3_1 _36007_ (.A(_13650_),
    .B(_12634_),
    .C(_13345_),
    .X(_13652_));
 sky130_fd_sc_hd__buf_6 _36008_ (.A(_13652_),
    .X(_13653_));
 sky130_fd_sc_hd__nor2_8 _36009_ (.A(_13651_),
    .B(_13653_),
    .Y(_13654_));
 sky130_fd_sc_hd__clkinv_4 _36010_ (.A(_13654_),
    .Y(_13655_));
 sky130_fd_sc_hd__buf_4 _36011_ (.A(_13655_),
    .X(_13656_));
 sky130_fd_sc_hd__a21o_1 _36012_ (.A1(_13646_),
    .A2(_13649_),
    .B1(_13656_),
    .X(_13657_));
 sky130_fd_sc_hd__a21oi_4 _36013_ (.A1(_13280_),
    .A2(_13281_),
    .B1(_13220_),
    .Y(_13658_));
 sky130_fd_sc_hd__a21oi_2 _36014_ (.A1(_13289_),
    .A2(_13282_),
    .B1(_13658_),
    .Y(_13659_));
 sky130_fd_sc_hd__nand3_2 _36015_ (.A(_13646_),
    .B(_13656_),
    .C(_13649_),
    .Y(_13660_));
 sky130_fd_sc_hd__nand3_4 _36016_ (.A(_13657_),
    .B(_13659_),
    .C(_13660_),
    .Y(_13661_));
 sky130_fd_sc_hd__a31oi_4 _36017_ (.A1(_13280_),
    .A2(_13281_),
    .A3(_13220_),
    .B1(_13284_),
    .Y(_13662_));
 sky130_fd_sc_hd__buf_4 _36018_ (.A(_13654_),
    .X(_13663_));
 sky130_fd_sc_hd__nand3_2 _36019_ (.A(_13646_),
    .B(_13649_),
    .C(_13663_),
    .Y(_13664_));
 sky130_fd_sc_hd__o2bb2ai_1 _36020_ (.A1_N(_13649_),
    .A2_N(_13646_),
    .B1(_13653_),
    .B2(_13651_),
    .Y(_13665_));
 sky130_fd_sc_hd__o211ai_4 _36021_ (.A1(_13658_),
    .A2(_13662_),
    .B1(_13664_),
    .C1(_13665_),
    .Y(_13666_));
 sky130_vsdinv _36022_ (.A(_13343_),
    .Y(_13667_));
 sky130_fd_sc_hd__and3_1 _36023_ (.A(_13337_),
    .B(_13348_),
    .C(_13349_),
    .X(_13668_));
 sky130_fd_sc_hd__or2_2 _36024_ (.A(_13667_),
    .B(_13668_),
    .X(_13669_));
 sky130_fd_sc_hd__a21oi_2 _36025_ (.A1(_13661_),
    .A2(_13666_),
    .B1(_13669_),
    .Y(_13670_));
 sky130_fd_sc_hd__nand3_2 _36026_ (.A(_13669_),
    .B(_13661_),
    .C(_13666_),
    .Y(_13671_));
 sky130_vsdinv _36027_ (.A(_13671_),
    .Y(_13672_));
 sky130_fd_sc_hd__o2bb2ai_2 _36028_ (.A1_N(_13614_),
    .A2_N(_13621_),
    .B1(_13670_),
    .B2(_13672_),
    .Y(_13673_));
 sky130_fd_sc_hd__a21bo_1 _36029_ (.A1(_13367_),
    .A2(_13293_),
    .B1_N(_13300_),
    .X(_13674_));
 sky130_fd_sc_hd__o21a_1 _36030_ (.A1(_13667_),
    .A2(_13668_),
    .B1(_13661_),
    .X(_13675_));
 sky130_fd_sc_hd__a21oi_2 _36031_ (.A1(_13675_),
    .A2(_13666_),
    .B1(_13670_),
    .Y(_13676_));
 sky130_fd_sc_hd__nand3_2 _36032_ (.A(_13621_),
    .B(_13614_),
    .C(_13676_),
    .Y(_13677_));
 sky130_fd_sc_hd__nand3_4 _36033_ (.A(_13673_),
    .B(_13674_),
    .C(_13677_),
    .Y(_13678_));
 sky130_fd_sc_hd__nand2_1 _36034_ (.A(_13661_),
    .B(_13666_),
    .Y(_13679_));
 sky130_fd_sc_hd__nor2_1 _36035_ (.A(_13667_),
    .B(_13668_),
    .Y(_13680_));
 sky130_fd_sc_hd__nand2_1 _36036_ (.A(_13679_),
    .B(_13680_),
    .Y(_13681_));
 sky130_fd_sc_hd__nand2_2 _36037_ (.A(_13681_),
    .B(_13671_),
    .Y(_13682_));
 sky130_fd_sc_hd__a21o_1 _36038_ (.A1(_13621_),
    .A2(_13614_),
    .B1(_13682_),
    .X(_13683_));
 sky130_fd_sc_hd__a21boi_4 _36039_ (.A1(_13367_),
    .A2(_13293_),
    .B1_N(_13300_),
    .Y(_13684_));
 sky130_fd_sc_hd__nand3_2 _36040_ (.A(_13621_),
    .B(_13614_),
    .C(_13682_),
    .Y(_13685_));
 sky130_fd_sc_hd__nand3_4 _36041_ (.A(_13683_),
    .B(_13684_),
    .C(_13685_),
    .Y(_13686_));
 sky130_fd_sc_hd__nand2_2 _36042_ (.A(_13348_),
    .B(_13650_),
    .Y(_13687_));
 sky130_vsdinv _36043_ (.A(_13687_),
    .Y(_13688_));
 sky130_fd_sc_hd__and2_2 _36044_ (.A(_13364_),
    .B(_13357_),
    .X(_13689_));
 sky130_fd_sc_hd__nor2_8 _36045_ (.A(_13688_),
    .B(_13689_),
    .Y(_13690_));
 sky130_fd_sc_hd__and3_1 _36046_ (.A(_13364_),
    .B(_13357_),
    .C(_13688_),
    .X(_13691_));
 sky130_fd_sc_hd__o2bb2ai_2 _36047_ (.A1_N(_13678_),
    .A2_N(_13686_),
    .B1(_13690_),
    .B2(_13691_),
    .Y(_13692_));
 sky130_fd_sc_hd__and3_1 _36048_ (.A(_13364_),
    .B(_13357_),
    .C(_13687_),
    .X(_13693_));
 sky130_fd_sc_hd__nor2_2 _36049_ (.A(_13687_),
    .B(_13689_),
    .Y(_13694_));
 sky130_fd_sc_hd__nor2_1 _36050_ (.A(_13693_),
    .B(_13694_),
    .Y(_13695_));
 sky130_vsdinv _36051_ (.A(_13695_),
    .Y(_13696_));
 sky130_fd_sc_hd__nand3_2 _36052_ (.A(_13686_),
    .B(_13678_),
    .C(_13696_),
    .Y(_13697_));
 sky130_fd_sc_hd__o21ai_2 _36053_ (.A1(_13382_),
    .A2(_13370_),
    .B1(_13381_),
    .Y(_13698_));
 sky130_fd_sc_hd__nand3_4 _36054_ (.A(_13692_),
    .B(_13697_),
    .C(_13698_),
    .Y(_13699_));
 sky130_fd_sc_hd__o2bb2ai_2 _36055_ (.A1_N(_13678_),
    .A2_N(_13686_),
    .B1(_13694_),
    .B2(_13693_),
    .Y(_13700_));
 sky130_fd_sc_hd__nand3_2 _36056_ (.A(_13686_),
    .B(_13678_),
    .C(_13695_),
    .Y(_13701_));
 sky130_fd_sc_hd__o21a_1 _36057_ (.A1(_13382_),
    .A2(_13370_),
    .B1(_13381_),
    .X(_13702_));
 sky130_fd_sc_hd__nand3_4 _36058_ (.A(_13700_),
    .B(_13701_),
    .C(_13702_),
    .Y(_13703_));
 sky130_fd_sc_hd__nand2_1 _36059_ (.A(_13699_),
    .B(_13703_),
    .Y(_13704_));
 sky130_fd_sc_hd__nand2_1 _36060_ (.A(_13704_),
    .B(_13385_),
    .Y(_13705_));
 sky130_fd_sc_hd__a21boi_2 _36061_ (.A1(_13384_),
    .A2(_13065_),
    .B1_N(_13390_),
    .Y(_13706_));
 sky130_fd_sc_hd__nand3b_2 _36062_ (.A_N(_13385_),
    .B(_13699_),
    .C(_13703_),
    .Y(_13707_));
 sky130_fd_sc_hd__nand3_4 _36063_ (.A(_13705_),
    .B(_13706_),
    .C(_13707_),
    .Y(_13708_));
 sky130_fd_sc_hd__o2bb2ai_2 _36064_ (.A1_N(_13699_),
    .A2_N(_13703_),
    .B1(_13090_),
    .B2(_13088_),
    .Y(_13709_));
 sky130_fd_sc_hd__nand2_1 _36065_ (.A(_13384_),
    .B(_13065_),
    .Y(_13710_));
 sky130_fd_sc_hd__nand2_1 _36066_ (.A(_13710_),
    .B(_13390_),
    .Y(_13711_));
 sky130_fd_sc_hd__nand3_2 _36067_ (.A(_13699_),
    .B(_13703_),
    .C(_13385_),
    .Y(_13712_));
 sky130_fd_sc_hd__nand3_4 _36068_ (.A(_13709_),
    .B(_13711_),
    .C(_13712_),
    .Y(_13713_));
 sky130_fd_sc_hd__nand2_2 _36069_ (.A(_13708_),
    .B(_13713_),
    .Y(_13714_));
 sky130_fd_sc_hd__nand3_1 _36070_ (.A(_13404_),
    .B(_13397_),
    .C(_13406_),
    .Y(_13715_));
 sky130_fd_sc_hd__nand2_2 _36071_ (.A(_13715_),
    .B(_13400_),
    .Y(_13716_));
 sky130_fd_sc_hd__xor2_4 _36072_ (.A(_13714_),
    .B(_13716_),
    .X(_02658_));
 sky130_vsdinv _36073_ (.A(_13653_),
    .Y(_13717_));
 sky130_fd_sc_hd__nand2_2 _36074_ (.A(_13717_),
    .B(_13650_),
    .Y(_13718_));
 sky130_vsdinv _36075_ (.A(_13718_),
    .Y(_13719_));
 sky130_fd_sc_hd__buf_4 _36076_ (.A(_13719_),
    .X(_13720_));
 sky130_fd_sc_hd__o21a_2 _36077_ (.A1(_13680_),
    .A2(_13679_),
    .B1(_13666_),
    .X(_13721_));
 sky130_fd_sc_hd__nor2_8 _36078_ (.A(_13720_),
    .B(_13721_),
    .Y(_13722_));
 sky130_fd_sc_hd__and3_2 _36079_ (.A(_13671_),
    .B(_13666_),
    .C(_13720_),
    .X(_13723_));
 sky130_fd_sc_hd__o21ai_2 _36080_ (.A1(_13619_),
    .A2(_13601_),
    .B1(_13611_),
    .Y(_13724_));
 sky130_fd_sc_hd__o21ai_4 _36081_ (.A1(_13594_),
    .A2(_13573_),
    .B1(_13583_),
    .Y(_13725_));
 sky130_fd_sc_hd__nand2_2 _36082_ (.A(_10281_),
    .B(_06649_),
    .Y(_13726_));
 sky130_fd_sc_hd__nand2_2 _36083_ (.A(_19587_),
    .B(_06650_),
    .Y(_13727_));
 sky130_fd_sc_hd__nor2_4 _36084_ (.A(_13726_),
    .B(_13727_),
    .Y(_13728_));
 sky130_fd_sc_hd__nor2_8 _36085_ (.A(net468),
    .B(net440),
    .Y(_13729_));
 sky130_fd_sc_hd__nand2_4 _36086_ (.A(_13726_),
    .B(_13727_),
    .Y(_13730_));
 sky130_fd_sc_hd__nand3b_2 _36087_ (.A_N(_13728_),
    .B(_13729_),
    .C(_13730_),
    .Y(_13731_));
 sky130_vsdinv _36088_ (.A(_13731_),
    .Y(_13732_));
 sky130_fd_sc_hd__buf_2 _36089_ (.A(_13728_),
    .X(_13733_));
 sky130_fd_sc_hd__inv_2 _36090_ (.A(_13730_),
    .Y(_13734_));
 sky130_vsdinv _36091_ (.A(_13729_),
    .Y(_13735_));
 sky130_fd_sc_hd__o21a_1 _36092_ (.A1(_13733_),
    .A2(_13734_),
    .B1(_13735_),
    .X(_13736_));
 sky130_fd_sc_hd__clkbuf_4 _36093_ (.A(_10830_),
    .X(_13737_));
 sky130_fd_sc_hd__nand3_2 _36094_ (.A(_11292_),
    .B(_13737_),
    .C(_05797_),
    .Y(_13738_));
 sky130_fd_sc_hd__nor2_2 _36095_ (.A(_19908_),
    .B(_13738_),
    .Y(_13739_));
 sky130_fd_sc_hd__a22oi_4 _36096_ (.A1(_12779_),
    .A2(_05797_),
    .B1(_08189_),
    .B2(_11292_),
    .Y(_13740_));
 sky130_fd_sc_hd__nand2_2 _36097_ (.A(_10828_),
    .B(_05799_),
    .Y(_13741_));
 sky130_fd_sc_hd__o21ai_4 _36098_ (.A1(_13739_),
    .A2(_13740_),
    .B1(_13741_),
    .Y(_13742_));
 sky130_fd_sc_hd__nand2_1 _36099_ (.A(_12401_),
    .B(_06827_),
    .Y(_13743_));
 sky130_fd_sc_hd__nand3b_4 _36100_ (.A_N(_13743_),
    .B(_13107_),
    .C(_08189_),
    .Y(_13744_));
 sky130_fd_sc_hd__buf_4 _36101_ (.A(_18474_),
    .X(_13745_));
 sky130_fd_sc_hd__o21ai_2 _36102_ (.A1(_19908_),
    .A2(_13745_),
    .B1(_13743_),
    .Y(_13746_));
 sky130_vsdinv _36103_ (.A(_13741_),
    .Y(_13747_));
 sky130_fd_sc_hd__nand3_4 _36104_ (.A(_13744_),
    .B(_13746_),
    .C(_13747_),
    .Y(_13748_));
 sky130_fd_sc_hd__o21ai_4 _36105_ (.A1(_13551_),
    .A2(_13550_),
    .B1(_13554_),
    .Y(_13749_));
 sky130_fd_sc_hd__a21oi_4 _36106_ (.A1(_13742_),
    .A2(_13748_),
    .B1(_13749_),
    .Y(_13750_));
 sky130_fd_sc_hd__o21ai_1 _36107_ (.A1(_19908_),
    .A2(_13738_),
    .B1(_13747_),
    .Y(_13751_));
 sky130_fd_sc_hd__o211a_4 _36108_ (.A1(_13740_),
    .A2(_13751_),
    .B1(_13749_),
    .C1(_13742_),
    .X(_13752_));
 sky130_fd_sc_hd__o22ai_4 _36109_ (.A1(_13732_),
    .A2(_13736_),
    .B1(_13750_),
    .B2(_13752_),
    .Y(_13753_));
 sky130_fd_sc_hd__o21ai_1 _36110_ (.A1(_13537_),
    .A2(_13542_),
    .B1(_13545_),
    .Y(_13754_));
 sky130_fd_sc_hd__o21ai_2 _36111_ (.A1(_13754_),
    .A2(_13558_),
    .B1(_13568_),
    .Y(_13755_));
 sky130_fd_sc_hd__nand2_1 _36112_ (.A(_13742_),
    .B(_13748_),
    .Y(_13756_));
 sky130_fd_sc_hd__a21oi_4 _36113_ (.A1(_13555_),
    .A2(_13556_),
    .B1(_13549_),
    .Y(_13757_));
 sky130_fd_sc_hd__nand2_4 _36114_ (.A(_13756_),
    .B(_13757_),
    .Y(_13758_));
 sky130_fd_sc_hd__nand3_4 _36115_ (.A(_13742_),
    .B(_13749_),
    .C(_13748_),
    .Y(_13759_));
 sky130_fd_sc_hd__nand3b_1 _36116_ (.A_N(_13728_),
    .B(_13735_),
    .C(_13730_),
    .Y(_13760_));
 sky130_fd_sc_hd__o21ai_1 _36117_ (.A1(_13733_),
    .A2(_13734_),
    .B1(_13729_),
    .Y(_13761_));
 sky130_fd_sc_hd__nand2_2 _36118_ (.A(_13760_),
    .B(_13761_),
    .Y(_13762_));
 sky130_fd_sc_hd__nand3_4 _36119_ (.A(_13758_),
    .B(_13759_),
    .C(_13762_),
    .Y(_13763_));
 sky130_fd_sc_hd__nand3_4 _36120_ (.A(_13753_),
    .B(_13755_),
    .C(_13763_),
    .Y(_13764_));
 sky130_fd_sc_hd__o21a_1 _36121_ (.A1(_13733_),
    .A2(_13734_),
    .B1(_13729_),
    .X(_13765_));
 sky130_fd_sc_hd__nor3_4 _36122_ (.A(_13733_),
    .B(_13729_),
    .C(_13734_),
    .Y(_13766_));
 sky130_fd_sc_hd__o22ai_4 _36123_ (.A1(_13765_),
    .A2(_13766_),
    .B1(_13750_),
    .B2(_13752_),
    .Y(_13767_));
 sky130_fd_sc_hd__a21oi_4 _36124_ (.A1(_13566_),
    .A2(_13567_),
    .B1(_13560_),
    .Y(_13768_));
 sky130_fd_sc_hd__o21ai_1 _36125_ (.A1(_13733_),
    .A2(_13734_),
    .B1(_13735_),
    .Y(_13769_));
 sky130_fd_sc_hd__nand2_2 _36126_ (.A(_13769_),
    .B(_13731_),
    .Y(_13770_));
 sky130_fd_sc_hd__nand3_4 _36127_ (.A(_13758_),
    .B(_13759_),
    .C(_13770_),
    .Y(_13771_));
 sky130_fd_sc_hd__nand3_4 _36128_ (.A(_13767_),
    .B(_13768_),
    .C(_13771_),
    .Y(_13772_));
 sky130_fd_sc_hd__nand2_2 _36129_ (.A(_10261_),
    .B(_06641_),
    .Y(_13773_));
 sky130_fd_sc_hd__nand3_2 _36130_ (.A(_13773_),
    .B(_13514_),
    .C(_11848_),
    .Y(_13774_));
 sky130_fd_sc_hd__nand2_2 _36131_ (.A(_19596_),
    .B(_06267_),
    .Y(_13775_));
 sky130_fd_sc_hd__nand3_2 _36132_ (.A(_13775_),
    .B(_11379_),
    .C(_07060_),
    .Y(_13776_));
 sky130_fd_sc_hd__o211ai_4 _36133_ (.A1(_08579_),
    .A2(_10993_),
    .B1(_13774_),
    .C1(_13776_),
    .Y(_13777_));
 sky130_fd_sc_hd__nand3b_4 _36134_ (.A_N(_13775_),
    .B(_08947_),
    .C(_06635_),
    .Y(_13778_));
 sky130_fd_sc_hd__nor2_2 _36135_ (.A(_08578_),
    .B(_10993_),
    .Y(_13779_));
 sky130_fd_sc_hd__nand2_1 _36136_ (.A(_13775_),
    .B(_13773_),
    .Y(_13780_));
 sky130_fd_sc_hd__nand3_4 _36137_ (.A(_13778_),
    .B(_13779_),
    .C(_13780_),
    .Y(_13781_));
 sky130_fd_sc_hd__nor2_2 _36138_ (.A(_13541_),
    .B(_13544_),
    .Y(_13782_));
 sky130_fd_sc_hd__o2bb2ai_4 _36139_ (.A1_N(_13777_),
    .A2_N(_13781_),
    .B1(_13537_),
    .B2(_13782_),
    .Y(_13783_));
 sky130_fd_sc_hd__o21ai_4 _36140_ (.A1(_13540_),
    .A2(_13536_),
    .B1(_13539_),
    .Y(_13784_));
 sky130_fd_sc_hd__nand3_4 _36141_ (.A(_13781_),
    .B(_13784_),
    .C(_13777_),
    .Y(_13785_));
 sky130_fd_sc_hd__a21oi_4 _36142_ (.A1(_13520_),
    .A2(_13518_),
    .B1(_13523_),
    .Y(_13786_));
 sky130_vsdinv _36143_ (.A(_13786_),
    .Y(_13787_));
 sky130_fd_sc_hd__a21oi_4 _36144_ (.A1(_13783_),
    .A2(_13785_),
    .B1(_13787_),
    .Y(_13788_));
 sky130_fd_sc_hd__and3_2 _36145_ (.A(_13783_),
    .B(_13785_),
    .C(_13787_),
    .X(_13789_));
 sky130_fd_sc_hd__o2bb2ai_2 _36146_ (.A1_N(_13764_),
    .A2_N(_13772_),
    .B1(_13788_),
    .B2(_13789_),
    .Y(_13790_));
 sky130_fd_sc_hd__nor2_8 _36147_ (.A(_13788_),
    .B(_13789_),
    .Y(_13791_));
 sky130_fd_sc_hd__nand3_4 _36148_ (.A(_13791_),
    .B(_13772_),
    .C(_13764_),
    .Y(_13792_));
 sky130_fd_sc_hd__nand3_4 _36149_ (.A(_13725_),
    .B(_13790_),
    .C(_13792_),
    .Y(_13793_));
 sky130_fd_sc_hd__a21oi_2 _36150_ (.A1(_13772_),
    .A2(_13764_),
    .B1(_13791_),
    .Y(_13794_));
 sky130_fd_sc_hd__a21oi_1 _36151_ (.A1(_13783_),
    .A2(_13785_),
    .B1(_13786_),
    .Y(_13795_));
 sky130_fd_sc_hd__a21oi_4 _36152_ (.A1(_13781_),
    .A2(_13777_),
    .B1(_13784_),
    .Y(_13796_));
 sky130_fd_sc_hd__nand2_2 _36153_ (.A(_13785_),
    .B(_13786_),
    .Y(_13797_));
 sky130_fd_sc_hd__nor2_1 _36154_ (.A(_13796_),
    .B(_13797_),
    .Y(_13798_));
 sky130_fd_sc_hd__o211a_1 _36155_ (.A1(_13795_),
    .A2(_13798_),
    .B1(_13764_),
    .C1(_13772_),
    .X(_13799_));
 sky130_fd_sc_hd__a21oi_4 _36156_ (.A1(_13577_),
    .A2(_13582_),
    .B1(_13575_),
    .Y(_13800_));
 sky130_fd_sc_hd__o21ai_4 _36157_ (.A1(_13794_),
    .A2(_13799_),
    .B1(_13800_),
    .Y(_13801_));
 sky130_fd_sc_hd__nand3_4 _36158_ (.A(_12468_),
    .B(_19612_),
    .C(_07051_),
    .Y(_13802_));
 sky130_fd_sc_hd__nor2_2 _36159_ (.A(_10732_),
    .B(_13802_),
    .Y(_13803_));
 sky130_fd_sc_hd__a22o_2 _36160_ (.A1(_19609_),
    .A2(_19879_),
    .B1(_19613_),
    .B2(_19875_),
    .X(_13804_));
 sky130_fd_sc_hd__nand2_2 _36161_ (.A(_19617_),
    .B(_08062_),
    .Y(_13805_));
 sky130_fd_sc_hd__nand3b_2 _36162_ (.A_N(_13803_),
    .B(_13804_),
    .C(_13805_),
    .Y(_13806_));
 sky130_fd_sc_hd__a21oi_2 _36163_ (.A1(_13478_),
    .A2(_13477_),
    .B1(_13475_),
    .Y(_13807_));
 sky130_fd_sc_hd__a22oi_4 _36164_ (.A1(_12468_),
    .A2(_19878_),
    .B1(_19612_),
    .B2(_07346_),
    .Y(_13808_));
 sky130_vsdinv _36165_ (.A(_13805_),
    .Y(_13809_));
 sky130_fd_sc_hd__o21ai_2 _36166_ (.A1(_13808_),
    .A2(_13803_),
    .B1(_13809_),
    .Y(_13810_));
 sky130_fd_sc_hd__nand3_4 _36167_ (.A(_13806_),
    .B(_13807_),
    .C(_13810_),
    .Y(_13811_));
 sky130_fd_sc_hd__nor2_2 _36168_ (.A(_13476_),
    .B(_13481_),
    .Y(_13812_));
 sky130_fd_sc_hd__o211ai_4 _36169_ (.A1(_10732_),
    .A2(_13802_),
    .B1(_13809_),
    .C1(_13804_),
    .Y(_13813_));
 sky130_fd_sc_hd__o21ai_2 _36170_ (.A1(_13808_),
    .A2(_13803_),
    .B1(_13805_),
    .Y(_13814_));
 sky130_fd_sc_hd__o211ai_4 _36171_ (.A1(_13475_),
    .A2(_13812_),
    .B1(_13813_),
    .C1(_13814_),
    .Y(_13815_));
 sky130_fd_sc_hd__a22oi_4 _36172_ (.A1(_11847_),
    .A2(_10149_),
    .B1(_11849_),
    .B2(_19866_),
    .Y(_13816_));
 sky130_fd_sc_hd__and4_1 _36173_ (.A(_07757_),
    .B(_19625_),
    .C(_08056_),
    .D(_19868_),
    .X(_13817_));
 sky130_fd_sc_hd__nand2_2 _36174_ (.A(_19627_),
    .B(_19862_),
    .Y(_13818_));
 sky130_vsdinv _36175_ (.A(_13818_),
    .Y(_13819_));
 sky130_fd_sc_hd__o21ai_2 _36176_ (.A1(_13816_),
    .A2(_13817_),
    .B1(_13819_),
    .Y(_13820_));
 sky130_fd_sc_hd__nand2_1 _36177_ (.A(_07484_),
    .B(_07701_),
    .Y(_13821_));
 sky130_fd_sc_hd__nand3b_4 _36178_ (.A_N(_13821_),
    .B(_19626_),
    .C(_10745_),
    .Y(_13822_));
 sky130_fd_sc_hd__a22o_1 _36179_ (.A1(_07934_),
    .A2(_07701_),
    .B1(_07825_),
    .B2(_09772_),
    .X(_13823_));
 sky130_fd_sc_hd__nand3_2 _36180_ (.A(_13822_),
    .B(_13818_),
    .C(_13823_),
    .Y(_13824_));
 sky130_fd_sc_hd__nand2_4 _36181_ (.A(_13820_),
    .B(_13824_),
    .Y(_13825_));
 sky130_fd_sc_hd__a21o_2 _36182_ (.A1(_13811_),
    .A2(_13815_),
    .B1(_13825_),
    .X(_13826_));
 sky130_fd_sc_hd__nand3_4 _36183_ (.A(_13811_),
    .B(_13815_),
    .C(_13825_),
    .Y(_13827_));
 sky130_fd_sc_hd__nand2_1 _36184_ (.A(_13530_),
    .B(_13532_),
    .Y(_13828_));
 sky130_fd_sc_hd__nand2_4 _36185_ (.A(_13828_),
    .B(_13526_),
    .Y(_13829_));
 sky130_fd_sc_hd__a21oi_4 _36186_ (.A1(_13826_),
    .A2(_13827_),
    .B1(_13829_),
    .Y(_13830_));
 sky130_fd_sc_hd__and3_1 _36187_ (.A(_13829_),
    .B(_13826_),
    .C(_13827_),
    .X(_13831_));
 sky130_fd_sc_hd__nand2_1 _36188_ (.A(_13497_),
    .B(_13487_),
    .Y(_13832_));
 sky130_fd_sc_hd__nand2_2 _36189_ (.A(_13832_),
    .B(_13483_),
    .Y(_13833_));
 sky130_vsdinv _36190_ (.A(_13833_),
    .Y(_13834_));
 sky130_fd_sc_hd__o21ai_1 _36191_ (.A1(_13830_),
    .A2(_13831_),
    .B1(_13834_),
    .Y(_13835_));
 sky130_vsdinv _36192_ (.A(_13835_),
    .Y(_13836_));
 sky130_fd_sc_hd__a21o_1 _36193_ (.A1(_13826_),
    .A2(_13827_),
    .B1(_13829_),
    .X(_13837_));
 sky130_fd_sc_hd__nand3_2 _36194_ (.A(_13829_),
    .B(_13826_),
    .C(_13827_),
    .Y(_13838_));
 sky130_fd_sc_hd__nand3_2 _36195_ (.A(_13837_),
    .B(_13838_),
    .C(_13833_),
    .Y(_13839_));
 sky130_vsdinv _36196_ (.A(_13839_),
    .Y(_13840_));
 sky130_fd_sc_hd__o2bb2ai_4 _36197_ (.A1_N(_13793_),
    .A2_N(_13801_),
    .B1(_13836_),
    .B2(_13840_),
    .Y(_13841_));
 sky130_fd_sc_hd__o21ai_1 _36198_ (.A1(_13830_),
    .A2(_13831_),
    .B1(_13833_),
    .Y(_13842_));
 sky130_fd_sc_hd__nand3_1 _36199_ (.A(_13837_),
    .B(_13838_),
    .C(_13834_),
    .Y(_13843_));
 sky130_fd_sc_hd__nand2_2 _36200_ (.A(_13842_),
    .B(_13843_),
    .Y(_13844_));
 sky130_fd_sc_hd__nand3_4 _36201_ (.A(_13801_),
    .B(_13793_),
    .C(_13844_),
    .Y(_13845_));
 sky130_fd_sc_hd__o21ai_4 _36202_ (.A1(_13591_),
    .A2(_13587_),
    .B1(_13597_),
    .Y(_13846_));
 sky130_fd_sc_hd__a21oi_4 _36203_ (.A1(_13841_),
    .A2(_13845_),
    .B1(_13846_),
    .Y(_13847_));
 sky130_fd_sc_hd__a21o_1 _36204_ (.A1(_13502_),
    .A2(_13511_),
    .B1(_13508_),
    .X(_13848_));
 sky130_fd_sc_hd__nand3_1 _36205_ (.A(_13502_),
    .B(_13511_),
    .C(_13508_),
    .Y(_13849_));
 sky130_fd_sc_hd__nand2_1 _36206_ (.A(_13576_),
    .B(_13584_),
    .Y(_13850_));
 sky130_fd_sc_hd__and2_1 _36207_ (.A(_13585_),
    .B(_13139_),
    .X(_13851_));
 sky130_fd_sc_hd__a22oi_2 _36208_ (.A1(_13848_),
    .A2(_13849_),
    .B1(_13850_),
    .B2(_13851_),
    .Y(_13852_));
 sky130_fd_sc_hd__o211a_2 _36209_ (.A1(_13588_),
    .A2(_13852_),
    .B1(_13845_),
    .C1(_13841_),
    .X(_13853_));
 sky130_fd_sc_hd__nand2_1 _36210_ (.A(_13511_),
    .B(_13508_),
    .Y(_13854_));
 sky130_fd_sc_hd__buf_6 _36211_ (.A(_11537_),
    .X(_13855_));
 sky130_fd_sc_hd__nand2_2 _36212_ (.A(_19631_),
    .B(_09972_),
    .Y(_13856_));
 sky130_fd_sc_hd__a21o_1 _36213_ (.A1(_10991_),
    .A2(_19855_),
    .B1(_13856_),
    .X(_13857_));
 sky130_fd_sc_hd__nand2_1 _36214_ (.A(_08873_),
    .B(_08773_),
    .Y(_13858_));
 sky130_fd_sc_hd__a21o_1 _36215_ (.A1(_19633_),
    .A2(_13413_),
    .B1(_13858_),
    .X(_13859_));
 sky130_fd_sc_hd__o211ai_4 _36216_ (.A1(net444),
    .A2(_13855_),
    .B1(_13857_),
    .C1(_13859_),
    .Y(_13860_));
 sky130_fd_sc_hd__nand3b_4 _36217_ (.A_N(_13856_),
    .B(_19636_),
    .C(_10643_),
    .Y(_13861_));
 sky130_fd_sc_hd__nor2_2 _36218_ (.A(net441),
    .B(_11537_),
    .Y(_13862_));
 sky130_fd_sc_hd__nand2_1 _36219_ (.A(_13856_),
    .B(_13858_),
    .Y(_13863_));
 sky130_fd_sc_hd__nand3_4 _36220_ (.A(_13861_),
    .B(_13862_),
    .C(_13863_),
    .Y(_13864_));
 sky130_fd_sc_hd__nand2_1 _36221_ (.A(_13860_),
    .B(_13864_),
    .Y(_13865_));
 sky130_fd_sc_hd__o21ai_1 _36222_ (.A1(_13489_),
    .A2(_13490_),
    .B1(_13493_),
    .Y(_13866_));
 sky130_fd_sc_hd__nand2_1 _36223_ (.A(_13489_),
    .B(_13490_),
    .Y(_13867_));
 sky130_fd_sc_hd__nand2_1 _36224_ (.A(_13866_),
    .B(_13867_),
    .Y(_13868_));
 sky130_fd_sc_hd__nand2_2 _36225_ (.A(_13865_),
    .B(_13868_),
    .Y(_13869_));
 sky130_fd_sc_hd__and2_1 _36226_ (.A(_13866_),
    .B(_13867_),
    .X(_13870_));
 sky130_fd_sc_hd__nand3_4 _36227_ (.A(_13870_),
    .B(_13864_),
    .C(_13860_),
    .Y(_13871_));
 sky130_fd_sc_hd__nand2_1 _36228_ (.A(_13869_),
    .B(_13871_),
    .Y(_13872_));
 sky130_fd_sc_hd__nor2_2 _36229_ (.A(_13415_),
    .B(_13418_),
    .Y(_13873_));
 sky130_fd_sc_hd__nor2_4 _36230_ (.A(_13412_),
    .B(_13873_),
    .Y(_13874_));
 sky130_vsdinv _36231_ (.A(_13874_),
    .Y(_13875_));
 sky130_fd_sc_hd__nand2_1 _36232_ (.A(_13872_),
    .B(_13875_),
    .Y(_13876_));
 sky130_fd_sc_hd__a21boi_2 _36233_ (.A1(_13424_),
    .A2(_13427_),
    .B1_N(_13420_),
    .Y(_13877_));
 sky130_fd_sc_hd__nand3_2 _36234_ (.A(_13869_),
    .B(_13871_),
    .C(_13874_),
    .Y(_13878_));
 sky130_fd_sc_hd__nand3_4 _36235_ (.A(_13876_),
    .B(_13877_),
    .C(_13878_),
    .Y(_13879_));
 sky130_fd_sc_hd__nand2_1 _36236_ (.A(_13872_),
    .B(_13874_),
    .Y(_13880_));
 sky130_fd_sc_hd__nand2_1 _36237_ (.A(_13428_),
    .B(_13420_),
    .Y(_13881_));
 sky130_fd_sc_hd__nand3_2 _36238_ (.A(_13869_),
    .B(_13871_),
    .C(_13875_),
    .Y(_13882_));
 sky130_fd_sc_hd__nand3_4 _36239_ (.A(_13880_),
    .B(_13881_),
    .C(_13882_),
    .Y(_13883_));
 sky130_fd_sc_hd__nand2_4 _36240_ (.A(_06156_),
    .B(_19834_),
    .Y(_13884_));
 sky130_fd_sc_hd__nand2_4 _36241_ (.A(_05883_),
    .B(_10504_),
    .Y(_13885_));
 sky130_fd_sc_hd__nor2_4 _36242_ (.A(_13884_),
    .B(_13885_),
    .Y(_13886_));
 sky130_fd_sc_hd__and2_1 _36243_ (.A(_13884_),
    .B(_13885_),
    .X(_13887_));
 sky130_fd_sc_hd__nand2_4 _36244_ (.A(_05732_),
    .B(_11597_),
    .Y(_13888_));
 sky130_fd_sc_hd__o21ai_2 _36245_ (.A1(_13886_),
    .A2(_13887_),
    .B1(_13888_),
    .Y(_13889_));
 sky130_vsdinv _36246_ (.A(_13888_),
    .Y(_13890_));
 sky130_fd_sc_hd__nand2_1 _36247_ (.A(_13884_),
    .B(_13885_),
    .Y(_13891_));
 sky130_fd_sc_hd__nand3b_2 _36248_ (.A_N(_13886_),
    .B(_13890_),
    .C(_13891_),
    .Y(_13892_));
 sky130_fd_sc_hd__nand2_4 _36249_ (.A(_13889_),
    .B(_13892_),
    .Y(_13893_));
 sky130_fd_sc_hd__a22oi_4 _36250_ (.A1(_19645_),
    .A2(_19849_),
    .B1(_19648_),
    .B2(_13248_),
    .Y(_13894_));
 sky130_fd_sc_hd__nand2_2 _36251_ (.A(_06411_),
    .B(_09359_),
    .Y(_13895_));
 sky130_fd_sc_hd__nand2_4 _36252_ (.A(_06169_),
    .B(_09817_),
    .Y(_13896_));
 sky130_fd_sc_hd__nor2_4 _36253_ (.A(_13895_),
    .B(_13896_),
    .Y(_13897_));
 sky130_fd_sc_hd__nand2_2 _36254_ (.A(net478),
    .B(_19839_),
    .Y(_13898_));
 sky130_fd_sc_hd__o21ai_4 _36255_ (.A1(_13894_),
    .A2(_13897_),
    .B1(_13898_),
    .Y(_13899_));
 sky130_fd_sc_hd__buf_6 _36256_ (.A(_10496_),
    .X(_13900_));
 sky130_fd_sc_hd__nand3_2 _36257_ (.A(_19645_),
    .B(_19648_),
    .C(_19849_),
    .Y(_13901_));
 sky130_fd_sc_hd__nand2_4 _36258_ (.A(_13895_),
    .B(_13896_),
    .Y(_13902_));
 sky130_vsdinv _36259_ (.A(_13898_),
    .Y(_13903_));
 sky130_fd_sc_hd__o211ai_4 _36260_ (.A1(_13900_),
    .A2(_13901_),
    .B1(_13902_),
    .C1(_13903_),
    .Y(_13904_));
 sky130_fd_sc_hd__nand2_1 _36261_ (.A(_13899_),
    .B(_13904_),
    .Y(_13905_));
 sky130_fd_sc_hd__a21oi_1 _36262_ (.A1(_13437_),
    .A2(_13436_),
    .B1(_13434_),
    .Y(_13906_));
 sky130_fd_sc_hd__nand2_1 _36263_ (.A(_13905_),
    .B(_13906_),
    .Y(_13907_));
 sky130_fd_sc_hd__a21o_2 _36264_ (.A1(_13437_),
    .A2(_13436_),
    .B1(_13434_),
    .X(_13908_));
 sky130_fd_sc_hd__nand3_4 _36265_ (.A(_13908_),
    .B(_13899_),
    .C(_13904_),
    .Y(_13909_));
 sky130_fd_sc_hd__nand2_1 _36266_ (.A(_13907_),
    .B(_13909_),
    .Y(_13910_));
 sky130_fd_sc_hd__nor2_2 _36267_ (.A(_13893_),
    .B(_13910_),
    .Y(_13911_));
 sky130_fd_sc_hd__and2_1 _36268_ (.A(_13910_),
    .B(_13893_),
    .X(_13912_));
 sky130_fd_sc_hd__o2bb2ai_4 _36269_ (.A1_N(_13879_),
    .A2_N(_13883_),
    .B1(_13911_),
    .B2(_13912_),
    .Y(_13913_));
 sky130_vsdinv _36270_ (.A(_13893_),
    .Y(_13914_));
 sky130_fd_sc_hd__nand2_1 _36271_ (.A(_13910_),
    .B(_13914_),
    .Y(_13915_));
 sky130_fd_sc_hd__nand3_1 _36272_ (.A(_13907_),
    .B(_13909_),
    .C(_13893_),
    .Y(_13916_));
 sky130_fd_sc_hd__nand2_2 _36273_ (.A(_13915_),
    .B(_13916_),
    .Y(_13917_));
 sky130_fd_sc_hd__nand3_4 _36274_ (.A(_13883_),
    .B(_13879_),
    .C(_13917_),
    .Y(_13918_));
 sky130_fd_sc_hd__a22oi_4 _36275_ (.A1(_13502_),
    .A2(_13854_),
    .B1(_13913_),
    .B2(_13918_),
    .Y(_13919_));
 sky130_vsdinv _36276_ (.A(_13511_),
    .Y(_13920_));
 sky130_fd_sc_hd__o211a_1 _36277_ (.A1(_13920_),
    .A2(_13510_),
    .B1(_13918_),
    .C1(_13913_),
    .X(_13921_));
 sky130_fd_sc_hd__and2_2 _36278_ (.A(_13464_),
    .B(_13463_),
    .X(_13922_));
 sky130_fd_sc_hd__o21ai_2 _36279_ (.A1(_13919_),
    .A2(_13921_),
    .B1(_13922_),
    .Y(_13923_));
 sky130_fd_sc_hd__a21oi_1 _36280_ (.A1(_13496_),
    .A2(_13498_),
    .B1(_13503_),
    .Y(_13924_));
 sky130_fd_sc_hd__o21ai_2 _36281_ (.A1(_13508_),
    .A2(_13924_),
    .B1(_13511_),
    .Y(_13925_));
 sky130_fd_sc_hd__a21o_1 _36282_ (.A1(_13913_),
    .A2(_13918_),
    .B1(_13925_),
    .X(_13926_));
 sky130_fd_sc_hd__nand3_4 _36283_ (.A(_13913_),
    .B(_13925_),
    .C(_13918_),
    .Y(_13927_));
 sky130_fd_sc_hd__nand3b_2 _36284_ (.A_N(_13922_),
    .B(_13926_),
    .C(_13927_),
    .Y(_13928_));
 sky130_fd_sc_hd__nand2_4 _36285_ (.A(_13923_),
    .B(_13928_),
    .Y(_13929_));
 sky130_fd_sc_hd__o21ai_2 _36286_ (.A1(_13847_),
    .A2(_13853_),
    .B1(_13929_),
    .Y(_13930_));
 sky130_fd_sc_hd__a21o_2 _36287_ (.A1(_13841_),
    .A2(_13845_),
    .B1(_13846_),
    .X(_13931_));
 sky130_fd_sc_hd__nand3_4 _36288_ (.A(_13846_),
    .B(_13841_),
    .C(_13845_),
    .Y(_13932_));
 sky130_fd_sc_hd__nand3b_2 _36289_ (.A_N(_13929_),
    .B(_13931_),
    .C(_13932_),
    .Y(_13933_));
 sky130_fd_sc_hd__nand3_4 _36290_ (.A(_13724_),
    .B(_13930_),
    .C(_13933_),
    .Y(_13934_));
 sky130_fd_sc_hd__a21oi_4 _36291_ (.A1(_13610_),
    .A2(_13612_),
    .B1(_13604_),
    .Y(_13935_));
 sky130_fd_sc_hd__nand3_4 _36292_ (.A(_13931_),
    .B(_13932_),
    .C(_13929_),
    .Y(_13936_));
 sky130_fd_sc_hd__o21bai_4 _36293_ (.A1(_13847_),
    .A2(_13853_),
    .B1_N(_13929_),
    .Y(_13937_));
 sky130_fd_sc_hd__nand3_4 _36294_ (.A(_13935_),
    .B(_13936_),
    .C(_13937_),
    .Y(_13938_));
 sky130_vsdinv _36295_ (.A(_13651_),
    .Y(_13939_));
 sky130_fd_sc_hd__a22o_1 _36296_ (.A1(_06327_),
    .A2(_19839_),
    .B1(_06838_),
    .B2(_10598_),
    .X(_13940_));
 sky130_fd_sc_hd__a21oi_4 _36297_ (.A1(_13940_),
    .A2(_13449_),
    .B1(_13445_),
    .Y(_13941_));
 sky130_fd_sc_hd__o21ai_4 _36298_ (.A1(_05450_),
    .A2(_06216_),
    .B1(_12274_),
    .Y(_13942_));
 sky130_fd_sc_hd__and3_4 _36299_ (.A(_18467_),
    .B(_05439_),
    .C(_05403_),
    .X(_13943_));
 sky130_fd_sc_hd__o21ai_4 _36300_ (.A1(_13942_),
    .A2(_13943_),
    .B1(_13307_),
    .Y(_13944_));
 sky130_fd_sc_hd__nand3_4 _36301_ (.A(_12274_),
    .B(_19661_),
    .C(_05842_),
    .Y(_13945_));
 sky130_fd_sc_hd__nand3b_4 _36302_ (.A_N(_13942_),
    .B(_13306_),
    .C(_13945_),
    .Y(_13946_));
 sky130_fd_sc_hd__nand3_4 _36303_ (.A(_13941_),
    .B(_13944_),
    .C(_13946_),
    .Y(_13947_));
 sky130_fd_sc_hd__nand2_1 _36304_ (.A(net477),
    .B(_09946_),
    .Y(_13948_));
 sky130_fd_sc_hd__nand3b_2 _36305_ (.A_N(_13948_),
    .B(_06160_),
    .C(_19835_),
    .Y(_13949_));
 sky130_fd_sc_hd__o21ai_2 _36306_ (.A1(_13447_),
    .A2(_13444_),
    .B1(_13949_),
    .Y(_13950_));
 sky130_fd_sc_hd__o21ai_4 _36307_ (.A1(_13942_),
    .A2(_13943_),
    .B1(_13310_),
    .Y(_13951_));
 sky130_fd_sc_hd__o211a_4 _36308_ (.A1(_05450_),
    .A2(_06216_),
    .B1(_12274_),
    .C1(_05259_),
    .X(_13952_));
 sky130_fd_sc_hd__nand2_8 _36309_ (.A(_13952_),
    .B(_13945_),
    .Y(_13953_));
 sky130_fd_sc_hd__nand3_4 _36310_ (.A(_13950_),
    .B(_13951_),
    .C(_13953_),
    .Y(_13954_));
 sky130_fd_sc_hd__a21oi_4 _36311_ (.A1(_13628_),
    .A2(_13310_),
    .B1(_13623_),
    .Y(_13955_));
 sky130_fd_sc_hd__a21oi_2 _36312_ (.A1(_13947_),
    .A2(_13954_),
    .B1(_13955_),
    .Y(_13956_));
 sky130_fd_sc_hd__and3_1 _36313_ (.A(_13947_),
    .B(_13954_),
    .C(_13955_),
    .X(_13957_));
 sky130_fd_sc_hd__a21oi_4 _36314_ (.A1(_13455_),
    .A2(_13451_),
    .B1(_13443_),
    .Y(_13958_));
 sky130_fd_sc_hd__o21ai_4 _36315_ (.A1(_13956_),
    .A2(_13957_),
    .B1(_13958_),
    .Y(_13959_));
 sky130_fd_sc_hd__o22ai_4 _36316_ (.A1(_13453_),
    .A2(_13454_),
    .B1(_13458_),
    .B2(_13440_),
    .Y(_13960_));
 sky130_fd_sc_hd__nand3_4 _36317_ (.A(_13947_),
    .B(_13954_),
    .C(_13955_),
    .Y(_13961_));
 sky130_fd_sc_hd__a21o_1 _36318_ (.A1(_13947_),
    .A2(_13954_),
    .B1(_13955_),
    .X(_13962_));
 sky130_fd_sc_hd__nand3_4 _36319_ (.A(_13960_),
    .B(_13961_),
    .C(_13962_),
    .Y(_13963_));
 sky130_fd_sc_hd__nand2_2 _36320_ (.A(_13631_),
    .B(_13636_),
    .Y(_13964_));
 sky130_fd_sc_hd__nand2_4 _36321_ (.A(_13964_),
    .B(_13635_),
    .Y(_13965_));
 sky130_fd_sc_hd__a21oi_4 _36322_ (.A1(_13959_),
    .A2(_13963_),
    .B1(_13965_),
    .Y(_13966_));
 sky130_vsdinv _36323_ (.A(_13635_),
    .Y(_13967_));
 sky130_vsdinv _36324_ (.A(_13964_),
    .Y(_13968_));
 sky130_fd_sc_hd__o211a_1 _36325_ (.A1(_13967_),
    .A2(_13968_),
    .B1(_13963_),
    .C1(_13959_),
    .X(_13969_));
 sky130_fd_sc_hd__a21oi_2 _36326_ (.A1(_13637_),
    .A2(_13638_),
    .B1(_13640_),
    .Y(_13970_));
 sky130_fd_sc_hd__o21ai_4 _36327_ (.A1(_13643_),
    .A2(_13970_),
    .B1(_13642_),
    .Y(_13971_));
 sky130_fd_sc_hd__o21bai_4 _36328_ (.A1(_13966_),
    .A2(_13969_),
    .B1_N(_13971_),
    .Y(_13972_));
 sky130_fd_sc_hd__a21o_1 _36329_ (.A1(_13959_),
    .A2(_13963_),
    .B1(_13965_),
    .X(_13973_));
 sky130_fd_sc_hd__nand3_4 _36330_ (.A(_13959_),
    .B(_13963_),
    .C(_13965_),
    .Y(_13974_));
 sky130_fd_sc_hd__nand3_4 _36331_ (.A(_13973_),
    .B(_13974_),
    .C(_13971_),
    .Y(_13975_));
 sky130_fd_sc_hd__a22oi_2 _36332_ (.A1(_13717_),
    .A2(_13939_),
    .B1(_13972_),
    .B2(_13975_),
    .Y(_13976_));
 sky130_fd_sc_hd__nand2_1 _36333_ (.A(_13971_),
    .B(_13974_),
    .Y(_13977_));
 sky130_fd_sc_hd__buf_2 _36334_ (.A(_13654_),
    .X(_13978_));
 sky130_fd_sc_hd__buf_4 _36335_ (.A(_13978_),
    .X(_13979_));
 sky130_fd_sc_hd__o211a_1 _36336_ (.A1(_13966_),
    .A2(_13977_),
    .B1(_13979_),
    .C1(_13972_),
    .X(_13980_));
 sky130_vsdinv _36337_ (.A(_13464_),
    .Y(_13981_));
 sky130_fd_sc_hd__nand2_1 _36338_ (.A(_13461_),
    .B(_13465_),
    .Y(_13982_));
 sky130_fd_sc_hd__o22ai_4 _36339_ (.A1(_13981_),
    .A2(_13982_),
    .B1(_13468_),
    .B2(_13470_),
    .Y(_13983_));
 sky130_fd_sc_hd__o21bai_2 _36340_ (.A1(_13976_),
    .A2(_13980_),
    .B1_N(_13983_),
    .Y(_13984_));
 sky130_fd_sc_hd__a21o_1 _36341_ (.A1(_13972_),
    .A2(_13975_),
    .B1(_13979_),
    .X(_13985_));
 sky130_fd_sc_hd__nand3_4 _36342_ (.A(_13972_),
    .B(_13979_),
    .C(_13975_),
    .Y(_13986_));
 sky130_fd_sc_hd__nand3_4 _36343_ (.A(_13985_),
    .B(_13986_),
    .C(_13983_),
    .Y(_13987_));
 sky130_fd_sc_hd__buf_2 _36344_ (.A(_13654_),
    .X(_13988_));
 sky130_fd_sc_hd__buf_6 _36345_ (.A(_13988_),
    .X(_13989_));
 sky130_fd_sc_hd__a21bo_1 _36346_ (.A1(_13989_),
    .A2(_13649_),
    .B1_N(_13646_),
    .X(_13990_));
 sky130_fd_sc_hd__a21oi_4 _36347_ (.A1(_13984_),
    .A2(_13987_),
    .B1(_13990_),
    .Y(_13991_));
 sky130_fd_sc_hd__nand3_2 _36348_ (.A(_13984_),
    .B(_13987_),
    .C(_13990_),
    .Y(_13992_));
 sky130_vsdinv _36349_ (.A(_13992_),
    .Y(_13993_));
 sky130_fd_sc_hd__o2bb2ai_4 _36350_ (.A1_N(_13934_),
    .A2_N(_13938_),
    .B1(_13991_),
    .B2(_13993_),
    .Y(_13994_));
 sky130_fd_sc_hd__nand2_1 _36351_ (.A(_13985_),
    .B(_13986_),
    .Y(_13995_));
 sky130_vsdinv _36352_ (.A(_13983_),
    .Y(_13996_));
 sky130_fd_sc_hd__a21boi_2 _36353_ (.A1(_13995_),
    .A2(_13996_),
    .B1_N(_13990_),
    .Y(_13997_));
 sky130_fd_sc_hd__a21oi_4 _36354_ (.A1(_13997_),
    .A2(_13987_),
    .B1(_13991_),
    .Y(_13998_));
 sky130_fd_sc_hd__nand3_4 _36355_ (.A(_13938_),
    .B(_13934_),
    .C(_13998_),
    .Y(_13999_));
 sky130_fd_sc_hd__nand2_1 _36356_ (.A(_13621_),
    .B(_13676_),
    .Y(_14000_));
 sky130_fd_sc_hd__nand2_4 _36357_ (.A(_14000_),
    .B(_13614_),
    .Y(_14001_));
 sky130_fd_sc_hd__a21oi_4 _36358_ (.A1(_13994_),
    .A2(_13999_),
    .B1(_14001_),
    .Y(_14002_));
 sky130_fd_sc_hd__and3_1 _36359_ (.A(_13605_),
    .B(_13607_),
    .C(_13613_),
    .X(_14003_));
 sky130_fd_sc_hd__a31oi_1 _36360_ (.A1(_13616_),
    .A2(_13615_),
    .A3(_13620_),
    .B1(_13682_),
    .Y(_14004_));
 sky130_fd_sc_hd__o211a_2 _36361_ (.A1(_14003_),
    .A2(_14004_),
    .B1(_13999_),
    .C1(_13994_),
    .X(_14005_));
 sky130_fd_sc_hd__o22ai_4 _36362_ (.A1(_13722_),
    .A2(_13723_),
    .B1(_14002_),
    .B2(_14005_),
    .Y(_14006_));
 sky130_fd_sc_hd__nand2_1 _36363_ (.A(_13686_),
    .B(_13696_),
    .Y(_14007_));
 sky130_fd_sc_hd__nand2_2 _36364_ (.A(_14007_),
    .B(_13678_),
    .Y(_14008_));
 sky130_fd_sc_hd__a21o_2 _36365_ (.A1(_13994_),
    .A2(_13999_),
    .B1(_14001_),
    .X(_14009_));
 sky130_fd_sc_hd__nand3_4 _36366_ (.A(_14001_),
    .B(_13994_),
    .C(_13999_),
    .Y(_14010_));
 sky130_fd_sc_hd__nor2_4 _36367_ (.A(_13723_),
    .B(_13722_),
    .Y(_14011_));
 sky130_fd_sc_hd__nand3_4 _36368_ (.A(_14009_),
    .B(_14010_),
    .C(_14011_),
    .Y(_14012_));
 sky130_fd_sc_hd__nand3_4 _36369_ (.A(_14006_),
    .B(_14008_),
    .C(_14012_),
    .Y(_14013_));
 sky130_vsdinv _36370_ (.A(_14011_),
    .Y(_14014_));
 sky130_fd_sc_hd__o21bai_2 _36371_ (.A1(_14002_),
    .A2(_14005_),
    .B1_N(_14014_),
    .Y(_14015_));
 sky130_fd_sc_hd__a21boi_4 _36372_ (.A1(_13686_),
    .A2(_13696_),
    .B1_N(_13678_),
    .Y(_14016_));
 sky130_fd_sc_hd__nand3_2 _36373_ (.A(_14009_),
    .B(_14010_),
    .C(_14014_),
    .Y(_14017_));
 sky130_fd_sc_hd__nand3_4 _36374_ (.A(_14015_),
    .B(_14016_),
    .C(_14017_),
    .Y(_14018_));
 sky130_fd_sc_hd__o2bb2ai_2 _36375_ (.A1_N(_14013_),
    .A2_N(_14018_),
    .B1(_13688_),
    .B2(_13689_),
    .Y(_14019_));
 sky130_fd_sc_hd__nand3_4 _36376_ (.A(_14018_),
    .B(_14013_),
    .C(_13690_),
    .Y(_14020_));
 sky130_fd_sc_hd__nand2_1 _36377_ (.A(_13703_),
    .B(_13385_),
    .Y(_14021_));
 sky130_fd_sc_hd__nand2_2 _36378_ (.A(_14021_),
    .B(_13699_),
    .Y(_14022_));
 sky130_fd_sc_hd__a21o_1 _36379_ (.A1(_14019_),
    .A2(_14020_),
    .B1(_14022_),
    .X(_14023_));
 sky130_fd_sc_hd__nand3_4 _36380_ (.A(_14019_),
    .B(_14022_),
    .C(_14020_),
    .Y(_14024_));
 sky130_fd_sc_hd__and2_1 _36381_ (.A(_14023_),
    .B(_14024_),
    .X(_14025_));
 sky130_vsdinv _36382_ (.A(_14025_),
    .Y(_14026_));
 sky130_fd_sc_hd__o2111ai_4 _36383_ (.A1(_13391_),
    .A2(_13395_),
    .B1(_13713_),
    .C1(_13708_),
    .D1(_13400_),
    .Y(_14027_));
 sky130_fd_sc_hd__nor2_4 _36384_ (.A(_14027_),
    .B(_13403_),
    .Y(_14028_));
 sky130_fd_sc_hd__and4_4 _36385_ (.A(_14028_),
    .B(_12039_),
    .C(_12041_),
    .D(_12384_),
    .X(_14029_));
 sky130_fd_sc_hd__a21boi_1 _36386_ (.A1(_13396_),
    .A2(_13708_),
    .B1_N(_13713_),
    .Y(_14030_));
 sky130_fd_sc_hd__o21ai_2 _36387_ (.A1(_14027_),
    .A2(_13406_),
    .B1(_14030_),
    .Y(_14031_));
 sky130_fd_sc_hd__a21oi_4 _36388_ (.A1(_12745_),
    .A2(_14028_),
    .B1(_14031_),
    .Y(_14032_));
 sky130_fd_sc_hd__a21boi_4 _36389_ (.A1(net409),
    .A2(_14029_),
    .B1_N(_14032_),
    .Y(_14033_));
 sky130_fd_sc_hd__nor2_8 _36390_ (.A(_14026_),
    .B(_14033_),
    .Y(_14034_));
 sky130_fd_sc_hd__and2_2 _36391_ (.A(_14033_),
    .B(_14026_),
    .X(_14035_));
 sky130_fd_sc_hd__nor2_8 _36392_ (.A(_14034_),
    .B(_14035_),
    .Y(_02659_));
 sky130_fd_sc_hd__o21ai_4 _36393_ (.A1(_14014_),
    .A2(_14002_),
    .B1(_14010_),
    .Y(_14036_));
 sky130_fd_sc_hd__nand2_1 _36394_ (.A(_13610_),
    .B(_13612_),
    .Y(_14037_));
 sky130_fd_sc_hd__a22oi_4 _36395_ (.A1(_14037_),
    .A2(_13611_),
    .B1(_13937_),
    .B2(_13936_),
    .Y(_14038_));
 sky130_fd_sc_hd__a21oi_4 _36396_ (.A1(_13938_),
    .A2(_13998_),
    .B1(_14038_),
    .Y(_14039_));
 sky130_fd_sc_hd__nand2_2 _36397_ (.A(_13932_),
    .B(_13929_),
    .Y(_14040_));
 sky130_fd_sc_hd__nand2_1 _36398_ (.A(_13835_),
    .B(_13839_),
    .Y(_14041_));
 sky130_fd_sc_hd__a21oi_2 _36399_ (.A1(_13790_),
    .A2(_13792_),
    .B1(_13725_),
    .Y(_14042_));
 sky130_fd_sc_hd__o21ai_4 _36400_ (.A1(_14041_),
    .A2(_14042_),
    .B1(_13793_),
    .Y(_14043_));
 sky130_fd_sc_hd__and3_2 _36401_ (.A(_13753_),
    .B(_13755_),
    .C(_13763_),
    .X(_14044_));
 sky130_fd_sc_hd__nand2_1 _36402_ (.A(_13783_),
    .B(_13785_),
    .Y(_14045_));
 sky130_fd_sc_hd__a2bb2oi_2 _36403_ (.A1_N(_13796_),
    .A2_N(_13797_),
    .B1(_13787_),
    .B2(_14045_),
    .Y(_14046_));
 sky130_fd_sc_hd__a31oi_4 _36404_ (.A1(_13768_),
    .A2(_13767_),
    .A3(_13771_),
    .B1(_14046_),
    .Y(_14047_));
 sky130_fd_sc_hd__a21oi_4 _36405_ (.A1(_13758_),
    .A2(_13762_),
    .B1(_13752_),
    .Y(_14048_));
 sky130_fd_sc_hd__nand2_4 _36406_ (.A(net469),
    .B(_19894_),
    .Y(_14049_));
 sky130_fd_sc_hd__nand2_4 _36407_ (.A(_19587_),
    .B(_07072_),
    .Y(_14050_));
 sky130_fd_sc_hd__nor2_4 _36408_ (.A(_14049_),
    .B(_14050_),
    .Y(_14051_));
 sky130_fd_sc_hd__and2_1 _36409_ (.A(_14049_),
    .B(_14050_),
    .X(_14052_));
 sky130_fd_sc_hd__nand2_4 _36410_ (.A(_10251_),
    .B(_06640_),
    .Y(_14053_));
 sky130_vsdinv _36411_ (.A(_14053_),
    .Y(_14054_));
 sky130_fd_sc_hd__o21ai_1 _36412_ (.A1(_14051_),
    .A2(_14052_),
    .B1(_14054_),
    .Y(_14055_));
 sky130_vsdinv _36413_ (.A(_14055_),
    .Y(_14056_));
 sky130_vsdinv _36414_ (.A(_14051_),
    .Y(_14057_));
 sky130_fd_sc_hd__nand2_4 _36415_ (.A(_14049_),
    .B(_14050_),
    .Y(_14058_));
 sky130_fd_sc_hd__nand3_2 _36416_ (.A(_14057_),
    .B(_14058_),
    .C(_14053_),
    .Y(_14059_));
 sky130_vsdinv _36417_ (.A(_14059_),
    .Y(_14060_));
 sky130_fd_sc_hd__nand3_2 _36418_ (.A(_11292_),
    .B(_13737_),
    .C(_05799_),
    .Y(_14061_));
 sky130_fd_sc_hd__nor2_2 _36419_ (.A(_19905_),
    .B(_14061_),
    .Y(_14062_));
 sky130_fd_sc_hd__a22oi_4 _36420_ (.A1(_13737_),
    .A2(_05811_),
    .B1(_05802_),
    .B2(_12402_),
    .Y(_14063_));
 sky130_fd_sc_hd__nand2_2 _36421_ (.A(_10828_),
    .B(_06119_),
    .Y(_14064_));
 sky130_fd_sc_hd__o21ai_4 _36422_ (.A1(_14062_),
    .A2(_14063_),
    .B1(_14064_),
    .Y(_14065_));
 sky130_fd_sc_hd__nand2_1 _36423_ (.A(_11079_),
    .B(_19901_),
    .Y(_14066_));
 sky130_fd_sc_hd__nand3b_4 _36424_ (.A_N(_14066_),
    .B(_12781_),
    .C(_05803_),
    .Y(_14067_));
 sky130_fd_sc_hd__o21ai_2 _36425_ (.A1(_19905_),
    .A2(_13745_),
    .B1(_14066_),
    .Y(_14068_));
 sky130_vsdinv _36426_ (.A(_14064_),
    .Y(_14069_));
 sky130_fd_sc_hd__nand3_4 _36427_ (.A(_14067_),
    .B(_14068_),
    .C(_14069_),
    .Y(_14070_));
 sky130_fd_sc_hd__o21ai_4 _36428_ (.A1(_13741_),
    .A2(_13740_),
    .B1(_13744_),
    .Y(_14071_));
 sky130_fd_sc_hd__a21oi_4 _36429_ (.A1(_14065_),
    .A2(_14070_),
    .B1(_14071_),
    .Y(_14072_));
 sky130_fd_sc_hd__o21ai_1 _36430_ (.A1(_19905_),
    .A2(_14061_),
    .B1(_14069_),
    .Y(_14073_));
 sky130_fd_sc_hd__o211a_4 _36431_ (.A1(_14063_),
    .A2(_14073_),
    .B1(_14071_),
    .C1(_14065_),
    .X(_14074_));
 sky130_fd_sc_hd__o22ai_4 _36432_ (.A1(_14056_),
    .A2(_14060_),
    .B1(_14072_),
    .B2(_14074_),
    .Y(_14075_));
 sky130_fd_sc_hd__a21o_2 _36433_ (.A1(_14065_),
    .A2(_14070_),
    .B1(_14071_),
    .X(_14076_));
 sky130_fd_sc_hd__nand3_4 _36434_ (.A(_14065_),
    .B(_14071_),
    .C(_14070_),
    .Y(_14077_));
 sky130_fd_sc_hd__nand3_1 _36435_ (.A(_14057_),
    .B(_14058_),
    .C(_14054_),
    .Y(_14078_));
 sky130_fd_sc_hd__o21ai_1 _36436_ (.A1(_14051_),
    .A2(_14052_),
    .B1(_14053_),
    .Y(_14079_));
 sky130_fd_sc_hd__nand2_2 _36437_ (.A(_14078_),
    .B(_14079_),
    .Y(_14080_));
 sky130_fd_sc_hd__nand3_4 _36438_ (.A(_14076_),
    .B(_14077_),
    .C(_14080_),
    .Y(_14081_));
 sky130_fd_sc_hd__nand3_4 _36439_ (.A(_14048_),
    .B(_14075_),
    .C(_14081_),
    .Y(_14082_));
 sky130_fd_sc_hd__a31o_2 _36440_ (.A1(_13730_),
    .A2(_19592_),
    .A3(_19892_),
    .B1(_13728_),
    .X(_14083_));
 sky130_fd_sc_hd__buf_4 _36441_ (.A(_10261_),
    .X(_14084_));
 sky130_fd_sc_hd__nand2_1 _36442_ (.A(_09722_),
    .B(_06634_),
    .Y(_14085_));
 sky130_fd_sc_hd__a21o_1 _36443_ (.A1(_14084_),
    .A2(_06804_),
    .B1(_14085_),
    .X(_14086_));
 sky130_fd_sc_hd__clkbuf_4 _36444_ (.A(_09485_),
    .X(_14087_));
 sky130_fd_sc_hd__nand2_1 _36445_ (.A(_08947_),
    .B(_19881_),
    .Y(_14088_));
 sky130_fd_sc_hd__a21o_1 _36446_ (.A1(_14087_),
    .A2(_07060_),
    .B1(_14088_),
    .X(_14089_));
 sky130_fd_sc_hd__nand2_2 _36447_ (.A(_19603_),
    .B(_07051_),
    .Y(_14090_));
 sky130_fd_sc_hd__nand3_4 _36448_ (.A(_14086_),
    .B(_14089_),
    .C(_14090_),
    .Y(_14091_));
 sky130_fd_sc_hd__nand3b_4 _36449_ (.A_N(_14085_),
    .B(_11379_),
    .C(_06804_),
    .Y(_14092_));
 sky130_vsdinv _36450_ (.A(_14090_),
    .Y(_14093_));
 sky130_fd_sc_hd__nand2_1 _36451_ (.A(_14085_),
    .B(_14088_),
    .Y(_14094_));
 sky130_fd_sc_hd__nand3_4 _36452_ (.A(_14092_),
    .B(_14093_),
    .C(_14094_),
    .Y(_14095_));
 sky130_fd_sc_hd__nand3_4 _36453_ (.A(_14083_),
    .B(_14091_),
    .C(_14095_),
    .Y(_14096_));
 sky130_fd_sc_hd__o21a_2 _36454_ (.A1(_13775_),
    .A2(_13773_),
    .B1(_13781_),
    .X(_14097_));
 sky130_fd_sc_hd__a21oi_4 _36455_ (.A1(_14091_),
    .A2(_14095_),
    .B1(_14083_),
    .Y(_14098_));
 sky130_fd_sc_hd__nor2_2 _36456_ (.A(_14097_),
    .B(_14098_),
    .Y(_14099_));
 sky130_fd_sc_hd__nor2_1 _36457_ (.A(_13733_),
    .B(_13729_),
    .Y(_14100_));
 sky130_fd_sc_hd__o2bb2ai_2 _36458_ (.A1_N(_14091_),
    .A2_N(_14095_),
    .B1(_13734_),
    .B2(_14100_),
    .Y(_14101_));
 sky130_fd_sc_hd__nand2_2 _36459_ (.A(_13781_),
    .B(_13778_),
    .Y(_14102_));
 sky130_fd_sc_hd__a21oi_4 _36460_ (.A1(_14101_),
    .A2(_14096_),
    .B1(_14102_),
    .Y(_14103_));
 sky130_fd_sc_hd__a21oi_4 _36461_ (.A1(_14096_),
    .A2(_14099_),
    .B1(_14103_),
    .Y(_14104_));
 sky130_fd_sc_hd__and3_1 _36462_ (.A(_14057_),
    .B(_14058_),
    .C(_14054_),
    .X(_14105_));
 sky130_vsdinv _36463_ (.A(_14079_),
    .Y(_14106_));
 sky130_fd_sc_hd__o22ai_4 _36464_ (.A1(_14105_),
    .A2(_14106_),
    .B1(_14072_),
    .B2(_14074_),
    .Y(_14107_));
 sky130_fd_sc_hd__o21ai_2 _36465_ (.A1(_13770_),
    .A2(_13750_),
    .B1(_13759_),
    .Y(_14108_));
 sky130_fd_sc_hd__nand2_2 _36466_ (.A(_14059_),
    .B(_14055_),
    .Y(_14109_));
 sky130_fd_sc_hd__nand3_4 _36467_ (.A(_14076_),
    .B(_14077_),
    .C(_14109_),
    .Y(_14110_));
 sky130_fd_sc_hd__nand3_4 _36468_ (.A(_14107_),
    .B(_14108_),
    .C(_14110_),
    .Y(_14111_));
 sky130_fd_sc_hd__nand3_4 _36469_ (.A(_14082_),
    .B(_14104_),
    .C(_14111_),
    .Y(_14112_));
 sky130_fd_sc_hd__and3_1 _36470_ (.A(_14101_),
    .B(_14102_),
    .C(_14096_),
    .X(_14113_));
 sky130_fd_sc_hd__o2bb2ai_2 _36471_ (.A1_N(_14111_),
    .A2_N(_14082_),
    .B1(_14103_),
    .B2(_14113_),
    .Y(_14114_));
 sky130_fd_sc_hd__o211ai_4 _36472_ (.A1(_14044_),
    .A2(_14047_),
    .B1(_14112_),
    .C1(_14114_),
    .Y(_14115_));
 sky130_fd_sc_hd__a21o_1 _36473_ (.A1(_14096_),
    .A2(_14099_),
    .B1(_14103_),
    .X(_14116_));
 sky130_fd_sc_hd__a21o_1 _36474_ (.A1(_14082_),
    .A2(_14111_),
    .B1(_14116_),
    .X(_14117_));
 sky130_fd_sc_hd__a21boi_4 _36475_ (.A1(_13791_),
    .A2(_13772_),
    .B1_N(_13764_),
    .Y(_14118_));
 sky130_fd_sc_hd__nand3_2 _36476_ (.A(_14116_),
    .B(_14082_),
    .C(_14111_),
    .Y(_14119_));
 sky130_fd_sc_hd__nand3_4 _36477_ (.A(_14117_),
    .B(_14118_),
    .C(_14119_),
    .Y(_14120_));
 sky130_fd_sc_hd__o22ai_4 _36478_ (.A1(_10732_),
    .A2(_13802_),
    .B1(_13805_),
    .B2(_13808_),
    .Y(_14121_));
 sky130_fd_sc_hd__a22oi_4 _36479_ (.A1(_19608_),
    .A2(_10733_),
    .B1(_12466_),
    .B2(_10957_),
    .Y(_14122_));
 sky130_fd_sc_hd__nand3_4 _36480_ (.A(_08908_),
    .B(_08550_),
    .C(_08735_),
    .Y(_14123_));
 sky130_fd_sc_hd__nor2_4 _36481_ (.A(_10960_),
    .B(_14123_),
    .Y(_14124_));
 sky130_fd_sc_hd__nand2_2 _36482_ (.A(_12470_),
    .B(_10395_),
    .Y(_14125_));
 sky130_vsdinv _36483_ (.A(_14125_),
    .Y(_14126_));
 sky130_fd_sc_hd__o21ai_2 _36484_ (.A1(_14122_),
    .A2(_14124_),
    .B1(_14126_),
    .Y(_14127_));
 sky130_fd_sc_hd__a22o_2 _36485_ (.A1(_19608_),
    .A2(_10733_),
    .B1(_19612_),
    .B2(_10957_),
    .X(_14128_));
 sky130_fd_sc_hd__o211ai_4 _36486_ (.A1(_11694_),
    .A2(_14123_),
    .B1(_14125_),
    .C1(_14128_),
    .Y(_14129_));
 sky130_fd_sc_hd__nand3b_4 _36487_ (.A_N(_14121_),
    .B(_14127_),
    .C(_14129_),
    .Y(_14130_));
 sky130_fd_sc_hd__o21ai_2 _36488_ (.A1(_14122_),
    .A2(_14124_),
    .B1(_14125_),
    .Y(_14131_));
 sky130_fd_sc_hd__o211ai_2 _36489_ (.A1(_11694_),
    .A2(_14123_),
    .B1(_14126_),
    .C1(_14128_),
    .Y(_14132_));
 sky130_fd_sc_hd__nand3_4 _36490_ (.A(_14131_),
    .B(_14121_),
    .C(_14132_),
    .Y(_14133_));
 sky130_fd_sc_hd__a22oi_4 _36491_ (.A1(_19622_),
    .A2(_08336_),
    .B1(_08565_),
    .B2(_08332_),
    .Y(_14134_));
 sky130_fd_sc_hd__nand2_2 _36492_ (.A(_07757_),
    .B(_08056_),
    .Y(_14135_));
 sky130_fd_sc_hd__nand2_2 _36493_ (.A(_08567_),
    .B(_19862_),
    .Y(_14136_));
 sky130_fd_sc_hd__nor2_4 _36494_ (.A(_14135_),
    .B(_14136_),
    .Y(_14137_));
 sky130_fd_sc_hd__a211o_1 _36495_ (.A1(_13408_),
    .A2(_13413_),
    .B1(_14134_),
    .C1(_14137_),
    .X(_14138_));
 sky130_fd_sc_hd__nand2_2 _36496_ (.A(_10364_),
    .B(_10453_),
    .Y(_14139_));
 sky130_vsdinv _36497_ (.A(_14139_),
    .Y(_14140_));
 sky130_fd_sc_hd__o21ai_2 _36498_ (.A1(_14134_),
    .A2(_14137_),
    .B1(_14140_),
    .Y(_14141_));
 sky130_fd_sc_hd__nand2_4 _36499_ (.A(_14138_),
    .B(_14141_),
    .Y(_14142_));
 sky130_fd_sc_hd__a21oi_2 _36500_ (.A1(_14130_),
    .A2(_14133_),
    .B1(_14142_),
    .Y(_14143_));
 sky130_fd_sc_hd__o21a_1 _36501_ (.A1(_14134_),
    .A2(_14137_),
    .B1(_14140_),
    .X(_14144_));
 sky130_fd_sc_hd__nor3_1 _36502_ (.A(_14140_),
    .B(_14134_),
    .C(_14137_),
    .Y(_14145_));
 sky130_fd_sc_hd__o211a_1 _36503_ (.A1(_14144_),
    .A2(_14145_),
    .B1(_14133_),
    .C1(_14130_),
    .X(_14146_));
 sky130_fd_sc_hd__nand2_4 _36504_ (.A(_13797_),
    .B(_13783_),
    .Y(_14147_));
 sky130_fd_sc_hd__o21ai_4 _36505_ (.A1(_14143_),
    .A2(_14146_),
    .B1(_14147_),
    .Y(_14148_));
 sky130_fd_sc_hd__a21o_2 _36506_ (.A1(_14130_),
    .A2(_14133_),
    .B1(_14142_),
    .X(_14149_));
 sky130_fd_sc_hd__nand3_4 _36507_ (.A(_14142_),
    .B(_14130_),
    .C(_14133_),
    .Y(_14150_));
 sky130_fd_sc_hd__o21ai_2 _36508_ (.A1(_13786_),
    .A2(_13796_),
    .B1(_13785_),
    .Y(_14151_));
 sky130_fd_sc_hd__nand3_4 _36509_ (.A(_14149_),
    .B(_14150_),
    .C(_14151_),
    .Y(_14152_));
 sky130_fd_sc_hd__nand2_1 _36510_ (.A(_13811_),
    .B(_13825_),
    .Y(_14153_));
 sky130_fd_sc_hd__nand2_4 _36511_ (.A(_14153_),
    .B(_13815_),
    .Y(_14154_));
 sky130_fd_sc_hd__a21oi_4 _36512_ (.A1(_14148_),
    .A2(_14152_),
    .B1(_14154_),
    .Y(_14155_));
 sky130_fd_sc_hd__and3_1 _36513_ (.A(_14148_),
    .B(_14152_),
    .C(_14154_),
    .X(_14156_));
 sky130_fd_sc_hd__o2bb2ai_2 _36514_ (.A1_N(_14115_),
    .A2_N(_14120_),
    .B1(_14155_),
    .B2(_14156_),
    .Y(_14157_));
 sky130_fd_sc_hd__nand2_1 _36515_ (.A(_14149_),
    .B(_14150_),
    .Y(_14158_));
 sky130_fd_sc_hd__a21boi_2 _36516_ (.A1(_14158_),
    .A2(_14147_),
    .B1_N(_14154_),
    .Y(_14159_));
 sky130_fd_sc_hd__a21oi_4 _36517_ (.A1(_14152_),
    .A2(_14159_),
    .B1(_14155_),
    .Y(_14160_));
 sky130_fd_sc_hd__nand3_4 _36518_ (.A(_14120_),
    .B(_14115_),
    .C(_14160_),
    .Y(_14161_));
 sky130_fd_sc_hd__nand3_4 _36519_ (.A(_14043_),
    .B(_14157_),
    .C(_14161_),
    .Y(_14162_));
 sky130_fd_sc_hd__a21boi_4 _36520_ (.A1(_13801_),
    .A2(_13844_),
    .B1_N(_13793_),
    .Y(_14163_));
 sky130_fd_sc_hd__nand2_1 _36521_ (.A(_14120_),
    .B(_14115_),
    .Y(_14164_));
 sky130_fd_sc_hd__nand2_1 _36522_ (.A(_14164_),
    .B(_14160_),
    .Y(_14165_));
 sky130_fd_sc_hd__nand3b_2 _36523_ (.A_N(_14160_),
    .B(_14115_),
    .C(_14120_),
    .Y(_14166_));
 sky130_fd_sc_hd__nand3_4 _36524_ (.A(_14163_),
    .B(_14165_),
    .C(_14166_),
    .Y(_14167_));
 sky130_fd_sc_hd__a31oi_4 _36525_ (.A1(_13829_),
    .A2(_13826_),
    .A3(_13827_),
    .B1(_13833_),
    .Y(_14168_));
 sky130_fd_sc_hd__a22oi_4 _36526_ (.A1(_08615_),
    .A2(_19854_),
    .B1(_08616_),
    .B2(_09075_),
    .Y(_14169_));
 sky130_fd_sc_hd__nand3_4 _36527_ (.A(_08190_),
    .B(_19635_),
    .C(_09076_),
    .Y(_14170_));
 sky130_fd_sc_hd__nor2_8 _36528_ (.A(_11537_),
    .B(_14170_),
    .Y(_14171_));
 sky130_fd_sc_hd__nand2_2 _36529_ (.A(_19641_),
    .B(_09358_),
    .Y(_14172_));
 sky130_vsdinv _36530_ (.A(_14172_),
    .Y(_14173_));
 sky130_fd_sc_hd__o21ai_2 _36531_ (.A1(_14169_),
    .A2(_14171_),
    .B1(_14173_),
    .Y(_14174_));
 sky130_fd_sc_hd__a21oi_2 _36532_ (.A1(_13823_),
    .A2(_13819_),
    .B1(_13817_),
    .Y(_14175_));
 sky130_fd_sc_hd__a22o_2 _36533_ (.A1(_08615_),
    .A2(_08773_),
    .B1(_08873_),
    .B2(_08787_),
    .X(_14176_));
 sky130_fd_sc_hd__o211ai_2 _36534_ (.A1(_11545_),
    .A2(_14170_),
    .B1(_14172_),
    .C1(_14176_),
    .Y(_14177_));
 sky130_fd_sc_hd__nand3_4 _36535_ (.A(_14174_),
    .B(_14175_),
    .C(_14177_),
    .Y(_14178_));
 sky130_fd_sc_hd__buf_2 _36536_ (.A(_14178_),
    .X(_14179_));
 sky130_fd_sc_hd__o21ai_4 _36537_ (.A1(_14169_),
    .A2(_14171_),
    .B1(_14172_),
    .Y(_14180_));
 sky130_fd_sc_hd__o211ai_4 _36538_ (.A1(_11545_),
    .A2(_14170_),
    .B1(_14173_),
    .C1(_14176_),
    .Y(_14181_));
 sky130_fd_sc_hd__o21ai_4 _36539_ (.A1(_13818_),
    .A2(_13816_),
    .B1(_13822_),
    .Y(_14182_));
 sky130_fd_sc_hd__nand3_4 _36540_ (.A(_14180_),
    .B(_14181_),
    .C(_14182_),
    .Y(_14183_));
 sky130_fd_sc_hd__nand2_1 _36541_ (.A(_13864_),
    .B(_13861_),
    .Y(_14184_));
 sky130_fd_sc_hd__clkbuf_2 _36542_ (.A(_14184_),
    .X(_14185_));
 sky130_fd_sc_hd__a21oi_2 _36543_ (.A1(_14179_),
    .A2(_14183_),
    .B1(_14185_),
    .Y(_14186_));
 sky130_fd_sc_hd__and3_1 _36544_ (.A(_14179_),
    .B(_14183_),
    .C(_14185_),
    .X(_14187_));
 sky130_fd_sc_hd__a21boi_4 _36545_ (.A1(_13869_),
    .A2(_13875_),
    .B1_N(_13871_),
    .Y(_14188_));
 sky130_fd_sc_hd__o21ai_4 _36546_ (.A1(_14186_),
    .A2(_14187_),
    .B1(_14188_),
    .Y(_14189_));
 sky130_fd_sc_hd__a21oi_1 _36547_ (.A1(_13860_),
    .A2(_13864_),
    .B1(_13870_),
    .Y(_14190_));
 sky130_fd_sc_hd__o21ai_2 _36548_ (.A1(_13874_),
    .A2(_14190_),
    .B1(_13871_),
    .Y(_14191_));
 sky130_fd_sc_hd__a21o_1 _36549_ (.A1(_14179_),
    .A2(_14183_),
    .B1(_14185_),
    .X(_14192_));
 sky130_fd_sc_hd__nand3_2 _36550_ (.A(_14179_),
    .B(_14183_),
    .C(_14185_),
    .Y(_14193_));
 sky130_fd_sc_hd__nand3_4 _36551_ (.A(_14191_),
    .B(_14192_),
    .C(_14193_),
    .Y(_14194_));
 sky130_fd_sc_hd__a21oi_4 _36552_ (.A1(_13903_),
    .A2(_13902_),
    .B1(_13897_),
    .Y(_14195_));
 sky130_fd_sc_hd__a22oi_4 _36553_ (.A1(_06411_),
    .A2(_11178_),
    .B1(_06618_),
    .B2(_11179_),
    .Y(_14196_));
 sky130_fd_sc_hd__nand3_4 _36554_ (.A(_06896_),
    .B(_19647_),
    .C(_19843_),
    .Y(_14197_));
 sky130_fd_sc_hd__nor2_4 _36555_ (.A(_09804_),
    .B(_14197_),
    .Y(_14198_));
 sky130_fd_sc_hd__o22ai_4 _36556_ (.A1(net473),
    .A2(_11206_),
    .B1(_14196_),
    .B2(_14198_),
    .Y(_14199_));
 sky130_fd_sc_hd__a22o_2 _36557_ (.A1(_06896_),
    .A2(_09950_),
    .B1(_06422_),
    .B2(_10488_),
    .X(_14200_));
 sky130_fd_sc_hd__nor2_4 _36558_ (.A(_11721_),
    .B(_11205_),
    .Y(_14201_));
 sky130_fd_sc_hd__o211ai_4 _36559_ (.A1(_09805_),
    .A2(_14197_),
    .B1(_14200_),
    .C1(_14201_),
    .Y(_14202_));
 sky130_fd_sc_hd__nand2_2 _36560_ (.A(_14199_),
    .B(_14202_),
    .Y(_14203_));
 sky130_fd_sc_hd__nor2_4 _36561_ (.A(_14195_),
    .B(_14203_),
    .Y(_14204_));
 sky130_fd_sc_hd__nand2_2 _36562_ (.A(_14203_),
    .B(_14195_),
    .Y(_14205_));
 sky130_fd_sc_hd__nand2_8 _36563_ (.A(_11184_),
    .B(_06013_),
    .Y(_14206_));
 sky130_vsdinv _36564_ (.A(_14206_),
    .Y(_14207_));
 sky130_fd_sc_hd__a22oi_4 _36565_ (.A1(_10737_),
    .A2(_11199_),
    .B1(_05737_),
    .B2(_11597_),
    .Y(_14208_));
 sky130_fd_sc_hd__nand2_4 _36566_ (.A(_07893_),
    .B(_19829_),
    .Y(_14209_));
 sky130_fd_sc_hd__nand2_4 _36567_ (.A(_06019_),
    .B(_10613_),
    .Y(_14210_));
 sky130_fd_sc_hd__nor2_8 _36568_ (.A(_14209_),
    .B(_14210_),
    .Y(_14211_));
 sky130_fd_sc_hd__nor3_4 _36569_ (.A(_14207_),
    .B(_14208_),
    .C(_14211_),
    .Y(_14212_));
 sky130_fd_sc_hd__o21a_1 _36570_ (.A1(_14208_),
    .A2(_14211_),
    .B1(_14207_),
    .X(_14213_));
 sky130_fd_sc_hd__nor2_4 _36571_ (.A(_14212_),
    .B(_14213_),
    .Y(_14214_));
 sky130_fd_sc_hd__nand3b_2 _36572_ (.A_N(_14204_),
    .B(_14205_),
    .C(_14214_),
    .Y(_14215_));
 sky130_fd_sc_hd__a21o_1 _36573_ (.A1(_13903_),
    .A2(_13902_),
    .B1(_13897_),
    .X(_14216_));
 sky130_fd_sc_hd__a21oi_4 _36574_ (.A1(_14199_),
    .A2(_14202_),
    .B1(_14216_),
    .Y(_14217_));
 sky130_fd_sc_hd__buf_6 _36575_ (.A(_11596_),
    .X(_14218_));
 sky130_fd_sc_hd__a211o_1 _36576_ (.A1(_14218_),
    .A2(net456),
    .B1(_14208_),
    .C1(_14211_),
    .X(_14219_));
 sky130_fd_sc_hd__o21ai_1 _36577_ (.A1(_14208_),
    .A2(_14211_),
    .B1(_14207_),
    .Y(_14220_));
 sky130_fd_sc_hd__nand2_2 _36578_ (.A(_14219_),
    .B(_14220_),
    .Y(_14221_));
 sky130_fd_sc_hd__o21ai_2 _36579_ (.A1(_14217_),
    .A2(_14204_),
    .B1(_14221_),
    .Y(_14222_));
 sky130_fd_sc_hd__nand2_4 _36580_ (.A(_14215_),
    .B(_14222_),
    .Y(_14223_));
 sky130_fd_sc_hd__a21oi_4 _36581_ (.A1(_14189_),
    .A2(_14194_),
    .B1(_14223_),
    .Y(_14224_));
 sky130_vsdinv _36582_ (.A(_14202_),
    .Y(_14225_));
 sky130_fd_sc_hd__nand2_2 _36583_ (.A(_14216_),
    .B(_14199_),
    .Y(_14226_));
 sky130_fd_sc_hd__o211a_1 _36584_ (.A1(_14225_),
    .A2(_14226_),
    .B1(_14214_),
    .C1(_14205_),
    .X(_14227_));
 sky130_fd_sc_hd__o21a_1 _36585_ (.A1(_14217_),
    .A2(_14204_),
    .B1(_14221_),
    .X(_14228_));
 sky130_fd_sc_hd__o211a_2 _36586_ (.A1(_14227_),
    .A2(_14228_),
    .B1(_14194_),
    .C1(_14189_),
    .X(_14229_));
 sky130_fd_sc_hd__o22ai_4 _36587_ (.A1(_13830_),
    .A2(_14168_),
    .B1(_14224_),
    .B2(_14229_),
    .Y(_14230_));
 sky130_fd_sc_hd__nor2_4 _36588_ (.A(_13830_),
    .B(_14168_),
    .Y(_14231_));
 sky130_fd_sc_hd__nand2_1 _36589_ (.A(_14189_),
    .B(_14194_),
    .Y(_14232_));
 sky130_fd_sc_hd__nor2_1 _36590_ (.A(_14227_),
    .B(_14228_),
    .Y(_14233_));
 sky130_fd_sc_hd__nand2_2 _36591_ (.A(_14232_),
    .B(_14233_),
    .Y(_14234_));
 sky130_fd_sc_hd__nand3_4 _36592_ (.A(_14223_),
    .B(_14189_),
    .C(_14194_),
    .Y(_14235_));
 sky130_fd_sc_hd__nand3_4 _36593_ (.A(_14231_),
    .B(_14234_),
    .C(_14235_),
    .Y(_14236_));
 sky130_vsdinv _36594_ (.A(_13883_),
    .Y(_14237_));
 sky130_fd_sc_hd__a21o_2 _36595_ (.A1(_13879_),
    .A2(_13917_),
    .B1(_14237_),
    .X(_14238_));
 sky130_fd_sc_hd__and3_2 _36596_ (.A(_14230_),
    .B(_14236_),
    .C(_14238_),
    .X(_14239_));
 sky130_fd_sc_hd__a21oi_4 _36597_ (.A1(_14230_),
    .A2(_14236_),
    .B1(_14238_),
    .Y(_14240_));
 sky130_fd_sc_hd__o2bb2ai_4 _36598_ (.A1_N(_14162_),
    .A2_N(_14167_),
    .B1(_14239_),
    .B2(_14240_),
    .Y(_14241_));
 sky130_fd_sc_hd__nor2_4 _36599_ (.A(_14240_),
    .B(_14239_),
    .Y(_14242_));
 sky130_fd_sc_hd__nand3_4 _36600_ (.A(_14242_),
    .B(_14167_),
    .C(_14162_),
    .Y(_14243_));
 sky130_fd_sc_hd__a22oi_4 _36601_ (.A1(_14040_),
    .A2(_13931_),
    .B1(_14241_),
    .B2(_14243_),
    .Y(_14244_));
 sky130_fd_sc_hd__a21o_1 _36602_ (.A1(_14230_),
    .A2(_14236_),
    .B1(_14238_),
    .X(_14245_));
 sky130_fd_sc_hd__nand3_2 _36603_ (.A(_14230_),
    .B(_14236_),
    .C(_14238_),
    .Y(_14246_));
 sky130_fd_sc_hd__nand2_4 _36604_ (.A(_14245_),
    .B(_14246_),
    .Y(_14247_));
 sky130_fd_sc_hd__a21o_1 _36605_ (.A1(_14167_),
    .A2(_14162_),
    .B1(_14247_),
    .X(_14248_));
 sky130_fd_sc_hd__nand3_4 _36606_ (.A(_14167_),
    .B(_14247_),
    .C(_14162_),
    .Y(_14249_));
 sky130_fd_sc_hd__nand2_2 _36607_ (.A(_14040_),
    .B(_13931_),
    .Y(_14250_));
 sky130_fd_sc_hd__a21oi_4 _36608_ (.A1(_14248_),
    .A2(_14249_),
    .B1(_14250_),
    .Y(_14251_));
 sky130_fd_sc_hd__a21oi_4 _36609_ (.A1(_13884_),
    .A2(_13885_),
    .B1(_13888_),
    .Y(_14252_));
 sky130_fd_sc_hd__nor2_2 _36610_ (.A(_13886_),
    .B(_14252_),
    .Y(_14253_));
 sky130_fd_sc_hd__nand3_4 _36611_ (.A(_14253_),
    .B(_13944_),
    .C(_13946_),
    .Y(_14254_));
 sky130_fd_sc_hd__o211ai_4 _36612_ (.A1(_13886_),
    .A2(_14252_),
    .B1(_13953_),
    .C1(_13951_),
    .Y(_14255_));
 sky130_fd_sc_hd__or2_4 _36613_ (.A(_13943_),
    .B(_13952_),
    .X(_14256_));
 sky130_fd_sc_hd__buf_4 _36614_ (.A(_14256_),
    .X(_14257_));
 sky130_fd_sc_hd__a21o_2 _36615_ (.A1(_14254_),
    .A2(_14255_),
    .B1(_14257_),
    .X(_14258_));
 sky130_fd_sc_hd__nand3_4 _36616_ (.A(_14254_),
    .B(_14255_),
    .C(_14257_),
    .Y(_14259_));
 sky130_fd_sc_hd__a21oi_4 _36617_ (.A1(_13899_),
    .A2(_13904_),
    .B1(_13908_),
    .Y(_14260_));
 sky130_fd_sc_hd__o21ai_4 _36618_ (.A1(_13893_),
    .A2(_14260_),
    .B1(_13909_),
    .Y(_14261_));
 sky130_fd_sc_hd__a21oi_4 _36619_ (.A1(_14258_),
    .A2(_14259_),
    .B1(_14261_),
    .Y(_14262_));
 sky130_fd_sc_hd__and3_2 _36620_ (.A(_14253_),
    .B(_13944_),
    .C(_13946_),
    .X(_14263_));
 sky130_fd_sc_hd__nand2_1 _36621_ (.A(_14255_),
    .B(_14257_),
    .Y(_14264_));
 sky130_fd_sc_hd__o211a_1 _36622_ (.A1(_14263_),
    .A2(_14264_),
    .B1(_14258_),
    .C1(_14261_),
    .X(_14265_));
 sky130_vsdinv _36623_ (.A(_13954_),
    .Y(_14266_));
 sky130_fd_sc_hd__a21oi_4 _36624_ (.A1(_13947_),
    .A2(_13955_),
    .B1(_14266_),
    .Y(_14267_));
 sky130_fd_sc_hd__o21ai_4 _36625_ (.A1(_14262_),
    .A2(_14265_),
    .B1(_14267_),
    .Y(_14268_));
 sky130_fd_sc_hd__a21o_1 _36626_ (.A1(_14258_),
    .A2(_14259_),
    .B1(_14261_),
    .X(_14269_));
 sky130_fd_sc_hd__nand3_4 _36627_ (.A(_14261_),
    .B(_14259_),
    .C(_14258_),
    .Y(_14270_));
 sky130_vsdinv _36628_ (.A(_14267_),
    .Y(_14271_));
 sky130_fd_sc_hd__nand3_4 _36629_ (.A(_14269_),
    .B(_14270_),
    .C(_14271_),
    .Y(_14272_));
 sky130_fd_sc_hd__nand2_2 _36630_ (.A(_13974_),
    .B(_13963_),
    .Y(_14273_));
 sky130_fd_sc_hd__a21oi_4 _36631_ (.A1(_14268_),
    .A2(_14272_),
    .B1(_14273_),
    .Y(_14274_));
 sky130_vsdinv _36632_ (.A(_13963_),
    .Y(_14275_));
 sky130_fd_sc_hd__nand2_1 _36633_ (.A(_13962_),
    .B(_13961_),
    .Y(_14276_));
 sky130_fd_sc_hd__a21boi_1 _36634_ (.A1(_14276_),
    .A2(_13958_),
    .B1_N(_13965_),
    .Y(_14277_));
 sky130_fd_sc_hd__o211a_2 _36635_ (.A1(_14275_),
    .A2(_14277_),
    .B1(_14272_),
    .C1(_14268_),
    .X(_14278_));
 sky130_fd_sc_hd__o21ai_2 _36636_ (.A1(_14274_),
    .A2(_14278_),
    .B1(_13979_),
    .Y(_14279_));
 sky130_fd_sc_hd__nand2_1 _36637_ (.A(_13922_),
    .B(_13927_),
    .Y(_14280_));
 sky130_fd_sc_hd__nand2_2 _36638_ (.A(_14280_),
    .B(_13926_),
    .Y(_14281_));
 sky130_fd_sc_hd__a21o_1 _36639_ (.A1(_14268_),
    .A2(_14272_),
    .B1(_14273_),
    .X(_14282_));
 sky130_fd_sc_hd__clkbuf_4 _36640_ (.A(_13655_),
    .X(_14283_));
 sky130_fd_sc_hd__nand3_2 _36641_ (.A(_14273_),
    .B(_14268_),
    .C(_14272_),
    .Y(_14284_));
 sky130_fd_sc_hd__nand3_2 _36642_ (.A(_14282_),
    .B(_14283_),
    .C(_14284_),
    .Y(_14285_));
 sky130_fd_sc_hd__nand3_4 _36643_ (.A(_14279_),
    .B(_14281_),
    .C(_14285_),
    .Y(_14286_));
 sky130_fd_sc_hd__o22ai_4 _36644_ (.A1(_13653_),
    .A2(_13651_),
    .B1(_14274_),
    .B2(_14278_),
    .Y(_14287_));
 sky130_fd_sc_hd__o21ai_4 _36645_ (.A1(_13922_),
    .A2(_13919_),
    .B1(_13927_),
    .Y(_14288_));
 sky130_fd_sc_hd__nand3_2 _36646_ (.A(_14282_),
    .B(_13979_),
    .C(_14284_),
    .Y(_14289_));
 sky130_fd_sc_hd__nand3_4 _36647_ (.A(_14287_),
    .B(_14288_),
    .C(_14289_),
    .Y(_14290_));
 sky130_fd_sc_hd__nand2_1 _36648_ (.A(_14286_),
    .B(_14290_),
    .Y(_14291_));
 sky130_vsdinv _36649_ (.A(_13975_),
    .Y(_14292_));
 sky130_fd_sc_hd__a21oi_1 _36650_ (.A1(_13973_),
    .A2(_13974_),
    .B1(_13971_),
    .Y(_14293_));
 sky130_fd_sc_hd__nor2_1 _36651_ (.A(_13656_),
    .B(_14293_),
    .Y(_14294_));
 sky130_fd_sc_hd__nor2_1 _36652_ (.A(_14292_),
    .B(_14294_),
    .Y(_14295_));
 sky130_fd_sc_hd__nand2_1 _36653_ (.A(_14291_),
    .B(_14295_),
    .Y(_14296_));
 sky130_vsdinv _36654_ (.A(_14295_),
    .Y(_14297_));
 sky130_fd_sc_hd__nand3_4 _36655_ (.A(_14297_),
    .B(_14286_),
    .C(_14290_),
    .Y(_14298_));
 sky130_fd_sc_hd__nand2_4 _36656_ (.A(_14296_),
    .B(_14298_),
    .Y(_14299_));
 sky130_fd_sc_hd__o21bai_4 _36657_ (.A1(_14244_),
    .A2(_14251_),
    .B1_N(_14299_),
    .Y(_14300_));
 sky130_fd_sc_hd__nor2_2 _36658_ (.A(_13929_),
    .B(_13847_),
    .Y(_14301_));
 sky130_fd_sc_hd__o211ai_4 _36659_ (.A1(_13853_),
    .A2(_14301_),
    .B1(_14243_),
    .C1(_14241_),
    .Y(_14302_));
 sky130_fd_sc_hd__nand3_4 _36660_ (.A(_14250_),
    .B(_14248_),
    .C(_14249_),
    .Y(_14303_));
 sky130_fd_sc_hd__nand3_4 _36661_ (.A(_14302_),
    .B(_14299_),
    .C(_14303_),
    .Y(_14304_));
 sky130_fd_sc_hd__buf_6 _36662_ (.A(_13718_),
    .X(_14305_));
 sky130_fd_sc_hd__nand2_2 _36663_ (.A(_13992_),
    .B(_13987_),
    .Y(_14306_));
 sky130_fd_sc_hd__nor2_4 _36664_ (.A(_14305_),
    .B(_14306_),
    .Y(_14307_));
 sky130_fd_sc_hd__nand2_1 _36665_ (.A(_14306_),
    .B(_14305_),
    .Y(_14308_));
 sky130_fd_sc_hd__or2b_1 _36666_ (.A(_14307_),
    .B_N(_14308_),
    .X(_14309_));
 sky130_fd_sc_hd__a31oi_4 _36667_ (.A1(_14039_),
    .A2(_14300_),
    .A3(_14304_),
    .B1(_14309_),
    .Y(_14310_));
 sky130_fd_sc_hd__nand2_2 _36668_ (.A(_13938_),
    .B(_13998_),
    .Y(_14311_));
 sky130_fd_sc_hd__nand2_1 _36669_ (.A(_14311_),
    .B(_13934_),
    .Y(_14312_));
 sky130_fd_sc_hd__nand3b_2 _36670_ (.A_N(_14299_),
    .B(_14302_),
    .C(_14303_),
    .Y(_14313_));
 sky130_fd_sc_hd__o21ai_2 _36671_ (.A1(_14244_),
    .A2(_14251_),
    .B1(_14299_),
    .Y(_14314_));
 sky130_fd_sc_hd__nand3_4 _36672_ (.A(_14312_),
    .B(_14313_),
    .C(_14314_),
    .Y(_14315_));
 sky130_fd_sc_hd__nand2_2 _36673_ (.A(_14310_),
    .B(_14315_),
    .Y(_14316_));
 sky130_fd_sc_hd__nand3_4 _36674_ (.A(_14039_),
    .B(_14300_),
    .C(_14304_),
    .Y(_14317_));
 sky130_vsdinv _36675_ (.A(_14308_),
    .Y(_14318_));
 sky130_fd_sc_hd__buf_2 _36676_ (.A(_14318_),
    .X(_14319_));
 sky130_fd_sc_hd__o2bb2ai_2 _36677_ (.A1_N(_14317_),
    .A2_N(_14315_),
    .B1(_14319_),
    .B2(_14307_),
    .Y(_14320_));
 sky130_fd_sc_hd__nand3_4 _36678_ (.A(_14036_),
    .B(_14316_),
    .C(_14320_),
    .Y(_14321_));
 sky130_fd_sc_hd__nor2_4 _36679_ (.A(_14307_),
    .B(_14318_),
    .Y(_14322_));
 sky130_fd_sc_hd__a21oi_2 _36680_ (.A1(_14315_),
    .A2(_14317_),
    .B1(_14322_),
    .Y(_14323_));
 sky130_fd_sc_hd__a22oi_4 _36681_ (.A1(_14311_),
    .A2(_13934_),
    .B1(_14300_),
    .B2(_14304_),
    .Y(_14324_));
 sky130_fd_sc_hd__nand2_1 _36682_ (.A(_14317_),
    .B(_14322_),
    .Y(_14325_));
 sky130_fd_sc_hd__nor2_2 _36683_ (.A(_14324_),
    .B(_14325_),
    .Y(_14326_));
 sky130_fd_sc_hd__a21oi_4 _36684_ (.A1(_14009_),
    .A2(_14011_),
    .B1(_14005_),
    .Y(_14327_));
 sky130_fd_sc_hd__o21ai_4 _36685_ (.A1(_14323_),
    .A2(_14326_),
    .B1(_14327_),
    .Y(_14328_));
 sky130_fd_sc_hd__buf_6 _36686_ (.A(net411),
    .X(_14329_));
 sky130_fd_sc_hd__buf_6 _36687_ (.A(_14329_),
    .X(_14330_));
 sky130_fd_sc_hd__buf_8 _36688_ (.A(_14330_),
    .X(_14331_));
 sky130_fd_sc_hd__clkbuf_4 _36689_ (.A(_14331_),
    .X(_14332_));
 sky130_fd_sc_hd__o2bb2ai_2 _36690_ (.A1_N(_14321_),
    .A2_N(_14328_),
    .B1(_14332_),
    .B2(_13721_),
    .Y(_14333_));
 sky130_fd_sc_hd__nand3_2 _36691_ (.A(_14328_),
    .B(_13722_),
    .C(_14321_),
    .Y(_14334_));
 sky130_vsdinv _36692_ (.A(_14012_),
    .Y(_14335_));
 sky130_fd_sc_hd__nand2_1 _36693_ (.A(_14006_),
    .B(_14008_),
    .Y(_14336_));
 sky130_fd_sc_hd__o2bb2ai_2 _36694_ (.A1_N(_13690_),
    .A2_N(_14018_),
    .B1(_14335_),
    .B2(_14336_),
    .Y(_14337_));
 sky130_fd_sc_hd__a21o_1 _36695_ (.A1(_14333_),
    .A2(_14334_),
    .B1(_14337_),
    .X(_14338_));
 sky130_fd_sc_hd__nand3_2 _36696_ (.A(_14333_),
    .B(_14337_),
    .C(_14334_),
    .Y(_14339_));
 sky130_fd_sc_hd__and2_2 _36697_ (.A(_14338_),
    .B(_14339_),
    .X(_14340_));
 sky130_fd_sc_hd__o21ai_4 _36698_ (.A1(_14026_),
    .A2(_14033_),
    .B1(_14024_),
    .Y(_14341_));
 sky130_fd_sc_hd__xor2_4 _36699_ (.A(_14340_),
    .B(_14341_),
    .X(_02660_));
 sky130_vsdinv _36700_ (.A(_14194_),
    .Y(_14342_));
 sky130_fd_sc_hd__and2_1 _36701_ (.A(_14223_),
    .B(_14189_),
    .X(_14343_));
 sky130_fd_sc_hd__a31o_1 _36702_ (.A1(_14181_),
    .A2(_14182_),
    .A3(_14180_),
    .B1(_14185_),
    .X(_14344_));
 sky130_fd_sc_hd__nor2_2 _36703_ (.A(_14173_),
    .B(_14171_),
    .Y(_14345_));
 sky130_fd_sc_hd__nand2_1 _36704_ (.A(_14135_),
    .B(_14136_),
    .Y(_14346_));
 sky130_fd_sc_hd__o21ai_2 _36705_ (.A1(_14135_),
    .A2(_14136_),
    .B1(_14139_),
    .Y(_14347_));
 sky130_fd_sc_hd__nand2_1 _36706_ (.A(_07744_),
    .B(_08787_),
    .Y(_14348_));
 sky130_fd_sc_hd__nand2_1 _36707_ (.A(_06921_),
    .B(_09358_),
    .Y(_14349_));
 sky130_fd_sc_hd__or2_2 _36708_ (.A(_14348_),
    .B(_14349_),
    .X(_14350_));
 sky130_fd_sc_hd__nor2_2 _36709_ (.A(net441),
    .B(_10497_),
    .Y(_14351_));
 sky130_fd_sc_hd__nand2_1 _36710_ (.A(_14348_),
    .B(_14349_),
    .Y(_14352_));
 sky130_fd_sc_hd__nand3_4 _36711_ (.A(_14350_),
    .B(_14351_),
    .C(_14352_),
    .Y(_14353_));
 sky130_fd_sc_hd__a21o_1 _36712_ (.A1(_10999_),
    .A2(_09820_),
    .B1(_14348_),
    .X(_14354_));
 sky130_fd_sc_hd__a21o_1 _36713_ (.A1(_10998_),
    .A2(_09362_),
    .B1(_14349_),
    .X(_14355_));
 sky130_fd_sc_hd__o211ai_4 _36714_ (.A1(net444),
    .A2(_10497_),
    .B1(_14354_),
    .C1(_14355_),
    .Y(_14356_));
 sky130_fd_sc_hd__a22oi_4 _36715_ (.A1(_14346_),
    .A2(_14347_),
    .B1(_14353_),
    .B2(_14356_),
    .Y(_14357_));
 sky130_fd_sc_hd__nor2_1 _36716_ (.A(_14139_),
    .B(_14134_),
    .Y(_14358_));
 sky130_fd_sc_hd__o211a_1 _36717_ (.A1(_14137_),
    .A2(_14358_),
    .B1(_14356_),
    .C1(_14353_),
    .X(_14359_));
 sky130_fd_sc_hd__o22ai_4 _36718_ (.A1(_14169_),
    .A2(_14345_),
    .B1(_14357_),
    .B2(_14359_),
    .Y(_14360_));
 sky130_fd_sc_hd__and2_1 _36719_ (.A(_14347_),
    .B(_14346_),
    .X(_14361_));
 sky130_fd_sc_hd__a21o_1 _36720_ (.A1(_14353_),
    .A2(_14356_),
    .B1(_14361_),
    .X(_14362_));
 sky130_fd_sc_hd__nand3_4 _36721_ (.A(_14361_),
    .B(_14353_),
    .C(_14356_),
    .Y(_14363_));
 sky130_fd_sc_hd__a21oi_4 _36722_ (.A1(_14176_),
    .A2(_14173_),
    .B1(_14171_),
    .Y(_14364_));
 sky130_vsdinv _36723_ (.A(_14364_),
    .Y(_14365_));
 sky130_fd_sc_hd__nand3_4 _36724_ (.A(_14362_),
    .B(_14363_),
    .C(_14365_),
    .Y(_14366_));
 sky130_fd_sc_hd__a22oi_4 _36725_ (.A1(_14179_),
    .A2(_14344_),
    .B1(_14360_),
    .B2(_14366_),
    .Y(_14367_));
 sky130_vsdinv _36726_ (.A(_14183_),
    .Y(_14368_));
 sky130_fd_sc_hd__and2_1 _36727_ (.A(_14178_),
    .B(_14184_),
    .X(_14369_));
 sky130_fd_sc_hd__o211a_1 _36728_ (.A1(_14368_),
    .A2(_14369_),
    .B1(_14366_),
    .C1(_14360_),
    .X(_14370_));
 sky130_fd_sc_hd__nand2_4 _36729_ (.A(_06608_),
    .B(_19838_),
    .Y(_14371_));
 sky130_fd_sc_hd__a21o_1 _36730_ (.A1(_06907_),
    .A2(_10487_),
    .B1(_14371_),
    .X(_14372_));
 sky130_fd_sc_hd__nand2_2 _36731_ (.A(_06416_),
    .B(_09933_),
    .Y(_14373_));
 sky130_fd_sc_hd__a21o_1 _36732_ (.A1(_08597_),
    .A2(_09946_),
    .B1(_14373_),
    .X(_14374_));
 sky130_fd_sc_hd__o211ai_4 _36733_ (.A1(net473),
    .A2(_10597_),
    .B1(_14372_),
    .C1(_14374_),
    .Y(_14375_));
 sky130_fd_sc_hd__nand3b_2 _36734_ (.A_N(_14371_),
    .B(_06618_),
    .C(_12639_),
    .Y(_14376_));
 sky130_fd_sc_hd__nor2_4 _36735_ (.A(_11721_),
    .B(_10596_),
    .Y(_14377_));
 sky130_fd_sc_hd__nand2_4 _36736_ (.A(_14371_),
    .B(_14373_),
    .Y(_14378_));
 sky130_fd_sc_hd__nand3_4 _36737_ (.A(_14376_),
    .B(_14377_),
    .C(_14378_),
    .Y(_14379_));
 sky130_fd_sc_hd__nand2_2 _36738_ (.A(_14375_),
    .B(_14379_),
    .Y(_14380_));
 sky130_fd_sc_hd__a21oi_4 _36739_ (.A1(_14201_),
    .A2(_14200_),
    .B1(_14198_),
    .Y(_14381_));
 sky130_fd_sc_hd__nand2_1 _36740_ (.A(_14380_),
    .B(_14381_),
    .Y(_14382_));
 sky130_fd_sc_hd__nand3b_2 _36741_ (.A_N(_14381_),
    .B(_14375_),
    .C(_14379_),
    .Y(_14383_));
 sky130_fd_sc_hd__nand2_4 _36742_ (.A(_07893_),
    .B(_10613_),
    .Y(_14384_));
 sky130_fd_sc_hd__nand2_8 _36743_ (.A(_11184_),
    .B(_05882_),
    .Y(_14385_));
 sky130_fd_sc_hd__nor2_8 _36744_ (.A(_14384_),
    .B(_14385_),
    .Y(_14386_));
 sky130_fd_sc_hd__nand2_2 _36745_ (.A(_14384_),
    .B(_14385_),
    .Y(_14387_));
 sky130_vsdinv _36746_ (.A(_14387_),
    .Y(_14388_));
 sky130_fd_sc_hd__o21ai_2 _36747_ (.A1(_14386_),
    .A2(_14388_),
    .B1(_14207_),
    .Y(_14389_));
 sky130_fd_sc_hd__nand3b_4 _36748_ (.A_N(_14386_),
    .B(_14206_),
    .C(_14387_),
    .Y(_14390_));
 sky130_fd_sc_hd__nand2_1 _36749_ (.A(_14389_),
    .B(_14390_),
    .Y(_14391_));
 sky130_fd_sc_hd__a21o_1 _36750_ (.A1(_14382_),
    .A2(_14383_),
    .B1(_14391_),
    .X(_14392_));
 sky130_fd_sc_hd__a22oi_4 _36751_ (.A1(_14389_),
    .A2(_14390_),
    .B1(_14380_),
    .B2(_14381_),
    .Y(_14393_));
 sky130_fd_sc_hd__nand2_1 _36752_ (.A(_14393_),
    .B(_14383_),
    .Y(_14394_));
 sky130_fd_sc_hd__nand2_4 _36753_ (.A(_14392_),
    .B(_14394_),
    .Y(_14395_));
 sky130_fd_sc_hd__o21bai_2 _36754_ (.A1(_14367_),
    .A2(_14370_),
    .B1_N(_14395_),
    .Y(_14396_));
 sky130_fd_sc_hd__a21boi_4 _36755_ (.A1(_14148_),
    .A2(_14154_),
    .B1_N(_14152_),
    .Y(_14397_));
 sky130_fd_sc_hd__a21o_1 _36756_ (.A1(_14185_),
    .A2(_14179_),
    .B1(_14368_),
    .X(_14398_));
 sky130_fd_sc_hd__a21o_1 _36757_ (.A1(_14360_),
    .A2(_14366_),
    .B1(_14398_),
    .X(_14399_));
 sky130_fd_sc_hd__nand3_4 _36758_ (.A(_14398_),
    .B(_14360_),
    .C(_14366_),
    .Y(_14400_));
 sky130_fd_sc_hd__nand3_4 _36759_ (.A(_14399_),
    .B(_14395_),
    .C(_14400_),
    .Y(_14401_));
 sky130_fd_sc_hd__nand3_4 _36760_ (.A(_14396_),
    .B(_14397_),
    .C(_14401_),
    .Y(_14402_));
 sky130_fd_sc_hd__o21ai_2 _36761_ (.A1(_14367_),
    .A2(_14370_),
    .B1(_14395_),
    .Y(_14403_));
 sky130_fd_sc_hd__nand3b_4 _36762_ (.A_N(_14395_),
    .B(_14399_),
    .C(_14400_),
    .Y(_14404_));
 sky130_fd_sc_hd__nand3b_4 _36763_ (.A_N(_14397_),
    .B(_14403_),
    .C(_14404_),
    .Y(_14405_));
 sky130_fd_sc_hd__o211a_4 _36764_ (.A1(_14342_),
    .A2(_14343_),
    .B1(_14402_),
    .C1(_14405_),
    .X(_14406_));
 sky130_fd_sc_hd__a21o_2 _36765_ (.A1(_14189_),
    .A2(_14223_),
    .B1(_14342_),
    .X(_14407_));
 sky130_fd_sc_hd__a21oi_4 _36766_ (.A1(_14405_),
    .A2(_14402_),
    .B1(_14407_),
    .Y(_14408_));
 sky130_fd_sc_hd__nand2_1 _36767_ (.A(_14082_),
    .B(_14104_),
    .Y(_14409_));
 sky130_fd_sc_hd__nand2_2 _36768_ (.A(_14409_),
    .B(_14111_),
    .Y(_14410_));
 sky130_fd_sc_hd__nand3_2 _36769_ (.A(_12780_),
    .B(_19576_),
    .C(_05977_),
    .Y(_14411_));
 sky130_fd_sc_hd__nor2_2 _36770_ (.A(_19902_),
    .B(_14411_),
    .Y(_14412_));
 sky130_fd_sc_hd__a22oi_4 _36771_ (.A1(_12401_),
    .A2(_06119_),
    .B1(net446),
    .B2(_12402_),
    .Y(_14413_));
 sky130_fd_sc_hd__nand2_2 _36772_ (.A(net498),
    .B(_05962_),
    .Y(_14414_));
 sky130_fd_sc_hd__o21ai_4 _36773_ (.A1(_14412_),
    .A2(_14413_),
    .B1(_14414_),
    .Y(_14415_));
 sky130_fd_sc_hd__nand2_1 _36774_ (.A(_11079_),
    .B(_06440_),
    .Y(_14416_));
 sky130_fd_sc_hd__nand3b_4 _36775_ (.A_N(_14416_),
    .B(_12781_),
    .C(net442),
    .Y(_14417_));
 sky130_fd_sc_hd__o21ai_2 _36776_ (.A1(_05799_),
    .A2(_13099_),
    .B1(_14416_),
    .Y(_14418_));
 sky130_vsdinv _36777_ (.A(_14414_),
    .Y(_14419_));
 sky130_fd_sc_hd__nand3_4 _36778_ (.A(_14417_),
    .B(_14418_),
    .C(_14419_),
    .Y(_14420_));
 sky130_fd_sc_hd__o21ai_4 _36779_ (.A1(_14064_),
    .A2(_14063_),
    .B1(_14067_),
    .Y(_14421_));
 sky130_fd_sc_hd__a21oi_4 _36780_ (.A1(_14415_),
    .A2(_14420_),
    .B1(_14421_),
    .Y(_14422_));
 sky130_fd_sc_hd__o21ai_1 _36781_ (.A1(_19902_),
    .A2(_14411_),
    .B1(_14419_),
    .Y(_14423_));
 sky130_fd_sc_hd__o211a_2 _36782_ (.A1(_14413_),
    .A2(_14423_),
    .B1(_14421_),
    .C1(_14415_),
    .X(_14424_));
 sky130_fd_sc_hd__nand2_2 _36783_ (.A(_11348_),
    .B(_06465_),
    .Y(_14425_));
 sky130_fd_sc_hd__nand2_2 _36784_ (.A(_10046_),
    .B(_06464_),
    .Y(_14426_));
 sky130_fd_sc_hd__nor2_4 _36785_ (.A(_14425_),
    .B(_14426_),
    .Y(_14427_));
 sky130_fd_sc_hd__nand2_2 _36786_ (.A(_14425_),
    .B(_14426_),
    .Y(_14428_));
 sky130_vsdinv _36787_ (.A(_14428_),
    .Y(_14429_));
 sky130_fd_sc_hd__nor2_4 _36788_ (.A(net468),
    .B(_08007_),
    .Y(_14430_));
 sky130_vsdinv _36789_ (.A(_14430_),
    .Y(_14431_));
 sky130_fd_sc_hd__o21ai_2 _36790_ (.A1(_14427_),
    .A2(_14429_),
    .B1(_14431_),
    .Y(_14432_));
 sky130_vsdinv _36791_ (.A(_14427_),
    .Y(_14433_));
 sky130_fd_sc_hd__nand3_2 _36792_ (.A(_14433_),
    .B(_14430_),
    .C(_14428_),
    .Y(_14434_));
 sky130_fd_sc_hd__nand2_4 _36793_ (.A(_14432_),
    .B(_14434_),
    .Y(_14435_));
 sky130_fd_sc_hd__o21ai_2 _36794_ (.A1(_14422_),
    .A2(_14424_),
    .B1(_14435_),
    .Y(_14436_));
 sky130_fd_sc_hd__o21ai_4 _36795_ (.A1(_14080_),
    .A2(_14072_),
    .B1(_14077_),
    .Y(_14437_));
 sky130_fd_sc_hd__a21o_1 _36796_ (.A1(_14415_),
    .A2(_14420_),
    .B1(_14421_),
    .X(_14438_));
 sky130_fd_sc_hd__nand3_4 _36797_ (.A(_14415_),
    .B(_14421_),
    .C(_14420_),
    .Y(_14439_));
 sky130_fd_sc_hd__nand3b_4 _36798_ (.A_N(_14435_),
    .B(_14438_),
    .C(_14439_),
    .Y(_14440_));
 sky130_fd_sc_hd__nand3_4 _36799_ (.A(_14436_),
    .B(_14437_),
    .C(_14440_),
    .Y(_14441_));
 sky130_fd_sc_hd__a21oi_4 _36800_ (.A1(_14076_),
    .A2(_14109_),
    .B1(_14074_),
    .Y(_14442_));
 sky130_fd_sc_hd__o21a_1 _36801_ (.A1(_14427_),
    .A2(_14429_),
    .B1(_14430_),
    .X(_14443_));
 sky130_fd_sc_hd__and3_1 _36802_ (.A(_14431_),
    .B(_14433_),
    .C(_14428_),
    .X(_14444_));
 sky130_fd_sc_hd__o22ai_4 _36803_ (.A1(_14443_),
    .A2(_14444_),
    .B1(_14422_),
    .B2(_14424_),
    .Y(_14445_));
 sky130_fd_sc_hd__nand3_4 _36804_ (.A(_14438_),
    .B(_14439_),
    .C(_14435_),
    .Y(_14446_));
 sky130_fd_sc_hd__nand3_4 _36805_ (.A(_14442_),
    .B(_14445_),
    .C(_14446_),
    .Y(_14447_));
 sky130_fd_sc_hd__nand2_1 _36806_ (.A(_10260_),
    .B(_06799_),
    .Y(_14448_));
 sky130_fd_sc_hd__a21o_1 _36807_ (.A1(_11379_),
    .A2(_07051_),
    .B1(_14448_),
    .X(_14449_));
 sky130_fd_sc_hd__nand2_1 _36808_ (.A(_09723_),
    .B(_07343_),
    .Y(_14450_));
 sky130_fd_sc_hd__a21o_1 _36809_ (.A1(_19597_),
    .A2(_07055_),
    .B1(_14450_),
    .X(_14451_));
 sky130_fd_sc_hd__clkbuf_4 _36810_ (.A(_09607_),
    .X(_14452_));
 sky130_fd_sc_hd__nand2_1 _36811_ (.A(_19603_),
    .B(_14452_),
    .Y(_14453_));
 sky130_fd_sc_hd__nand3_4 _36812_ (.A(_14449_),
    .B(_14451_),
    .C(_14453_),
    .Y(_14454_));
 sky130_fd_sc_hd__nand3_2 _36813_ (.A(_19597_),
    .B(_08947_),
    .C(_07055_),
    .Y(_14455_));
 sky130_fd_sc_hd__nand2_1 _36814_ (.A(_14448_),
    .B(_14450_),
    .Y(_14456_));
 sky130_fd_sc_hd__o2111ai_4 _36815_ (.A1(_08447_),
    .A2(_14455_),
    .B1(_19603_),
    .C1(_14452_),
    .D1(_14456_),
    .Y(_14457_));
 sky130_fd_sc_hd__nand2_1 _36816_ (.A(_14454_),
    .B(_14457_),
    .Y(_14458_));
 sky130_fd_sc_hd__o21ai_4 _36817_ (.A1(_14049_),
    .A2(_14050_),
    .B1(_14053_),
    .Y(_14459_));
 sky130_fd_sc_hd__nand2_1 _36818_ (.A(_14459_),
    .B(_14058_),
    .Y(_14460_));
 sky130_fd_sc_hd__nand2_2 _36819_ (.A(_14458_),
    .B(_14460_),
    .Y(_14461_));
 sky130_fd_sc_hd__nand3b_4 _36820_ (.A_N(_14460_),
    .B(_14454_),
    .C(_14457_),
    .Y(_14462_));
 sky130_fd_sc_hd__nand2_4 _36821_ (.A(_14095_),
    .B(_14092_),
    .Y(_14463_));
 sky130_fd_sc_hd__a21oi_2 _36822_ (.A1(_14461_),
    .A2(_14462_),
    .B1(_14463_),
    .Y(_14464_));
 sky130_fd_sc_hd__a21oi_2 _36823_ (.A1(_14049_),
    .A2(_14050_),
    .B1(_14053_),
    .Y(_14465_));
 sky130_fd_sc_hd__o211a_2 _36824_ (.A1(_14051_),
    .A2(_14465_),
    .B1(_14457_),
    .C1(_14454_),
    .X(_14466_));
 sky130_fd_sc_hd__nand2_4 _36825_ (.A(_14461_),
    .B(_14463_),
    .Y(_14467_));
 sky130_fd_sc_hd__nor2_2 _36826_ (.A(_14466_),
    .B(_14467_),
    .Y(_14468_));
 sky130_fd_sc_hd__o2bb2ai_4 _36827_ (.A1_N(_14441_),
    .A2_N(_14447_),
    .B1(_14464_),
    .B2(_14468_),
    .Y(_14469_));
 sky130_fd_sc_hd__a22oi_4 _36828_ (.A1(_14058_),
    .A2(_14459_),
    .B1(_14454_),
    .B2(_14457_),
    .Y(_14470_));
 sky130_fd_sc_hd__o21bai_2 _36829_ (.A1(_14470_),
    .A2(_14466_),
    .B1_N(_14463_),
    .Y(_14471_));
 sky130_fd_sc_hd__o21ai_4 _36830_ (.A1(_14466_),
    .A2(_14467_),
    .B1(_14471_),
    .Y(_14472_));
 sky130_vsdinv _36831_ (.A(_14472_),
    .Y(_14473_));
 sky130_fd_sc_hd__nand3_4 _36832_ (.A(_14473_),
    .B(_14441_),
    .C(_14447_),
    .Y(_14474_));
 sky130_fd_sc_hd__nand3_4 _36833_ (.A(_14410_),
    .B(_14469_),
    .C(_14474_),
    .Y(_14475_));
 sky130_fd_sc_hd__nand2_1 _36834_ (.A(_14447_),
    .B(_14441_),
    .Y(_14476_));
 sky130_fd_sc_hd__nand2_1 _36835_ (.A(_14476_),
    .B(_14473_),
    .Y(_14477_));
 sky130_fd_sc_hd__a21boi_4 _36836_ (.A1(_14082_),
    .A2(_14104_),
    .B1_N(_14111_),
    .Y(_14478_));
 sky130_fd_sc_hd__nand3_2 _36837_ (.A(_14447_),
    .B(_14441_),
    .C(_14472_),
    .Y(_14479_));
 sky130_fd_sc_hd__nand3_4 _36838_ (.A(_14477_),
    .B(_14478_),
    .C(_14479_),
    .Y(_14480_));
 sky130_fd_sc_hd__nand2_4 _36839_ (.A(_08153_),
    .B(_19871_),
    .Y(_14481_));
 sky130_fd_sc_hd__nand2_4 _36840_ (.A(_08541_),
    .B(_07701_),
    .Y(_14482_));
 sky130_fd_sc_hd__nor2_8 _36841_ (.A(_14481_),
    .B(_14482_),
    .Y(_14483_));
 sky130_fd_sc_hd__and2_1 _36842_ (.A(_14481_),
    .B(_14482_),
    .X(_14484_));
 sky130_fd_sc_hd__nand2_2 _36843_ (.A(_12470_),
    .B(_09772_),
    .Y(_14485_));
 sky130_fd_sc_hd__o21ai_2 _36844_ (.A1(_14483_),
    .A2(_14484_),
    .B1(_14485_),
    .Y(_14486_));
 sky130_fd_sc_hd__a21o_1 _36845_ (.A1(_14128_),
    .A2(_14126_),
    .B1(_14124_),
    .X(_14487_));
 sky130_fd_sc_hd__nand2_2 _36846_ (.A(_14481_),
    .B(_14482_),
    .Y(_14488_));
 sky130_vsdinv _36847_ (.A(_14485_),
    .Y(_14489_));
 sky130_fd_sc_hd__nand3b_2 _36848_ (.A_N(_14483_),
    .B(_14488_),
    .C(_14489_),
    .Y(_14490_));
 sky130_fd_sc_hd__nand3_4 _36849_ (.A(_14486_),
    .B(_14487_),
    .C(_14490_),
    .Y(_14491_));
 sky130_fd_sc_hd__o21ai_2 _36850_ (.A1(_14483_),
    .A2(_14484_),
    .B1(_14489_),
    .Y(_14492_));
 sky130_fd_sc_hd__nand3b_2 _36851_ (.A_N(_14483_),
    .B(_14488_),
    .C(_14485_),
    .Y(_14493_));
 sky130_fd_sc_hd__a21oi_2 _36852_ (.A1(_14128_),
    .A2(_14126_),
    .B1(_14124_),
    .Y(_14494_));
 sky130_fd_sc_hd__nand3_4 _36853_ (.A(_14492_),
    .B(_14493_),
    .C(_14494_),
    .Y(_14495_));
 sky130_fd_sc_hd__nand2_1 _36854_ (.A(_19622_),
    .B(_08332_),
    .Y(_14496_));
 sky130_fd_sc_hd__nand2_2 _36855_ (.A(_08565_),
    .B(_10459_),
    .Y(_14497_));
 sky130_fd_sc_hd__nor2_2 _36856_ (.A(_14496_),
    .B(_14497_),
    .Y(_14498_));
 sky130_fd_sc_hd__nand2_1 _36857_ (.A(_14496_),
    .B(_14497_),
    .Y(_14499_));
 sky130_vsdinv _36858_ (.A(_14499_),
    .Y(_14500_));
 sky130_fd_sc_hd__clkbuf_4 _36859_ (.A(_11232_),
    .X(_14501_));
 sky130_fd_sc_hd__nand2_1 _36860_ (.A(_11003_),
    .B(_14501_),
    .Y(_14502_));
 sky130_fd_sc_hd__o21bai_1 _36861_ (.A1(_14498_),
    .A2(_14500_),
    .B1_N(_14502_),
    .Y(_14503_));
 sky130_fd_sc_hd__nand3b_2 _36862_ (.A_N(_14498_),
    .B(_14502_),
    .C(_14499_),
    .Y(_14504_));
 sky130_fd_sc_hd__nand2_2 _36863_ (.A(_14503_),
    .B(_14504_),
    .Y(_14505_));
 sky130_fd_sc_hd__a21o_1 _36864_ (.A1(_14491_),
    .A2(_14495_),
    .B1(_14505_),
    .X(_14506_));
 sky130_fd_sc_hd__nand3_4 _36865_ (.A(_14505_),
    .B(_14491_),
    .C(_14495_),
    .Y(_14507_));
 sky130_fd_sc_hd__o21ai_4 _36866_ (.A1(_14097_),
    .A2(_14098_),
    .B1(_14096_),
    .Y(_14508_));
 sky130_fd_sc_hd__a21o_2 _36867_ (.A1(_14506_),
    .A2(_14507_),
    .B1(_14508_),
    .X(_14509_));
 sky130_fd_sc_hd__nand3_4 _36868_ (.A(_14506_),
    .B(_14507_),
    .C(_14508_),
    .Y(_14510_));
 sky130_fd_sc_hd__nand2_4 _36869_ (.A(_14150_),
    .B(_14133_),
    .Y(_14511_));
 sky130_fd_sc_hd__a21oi_4 _36870_ (.A1(_14509_),
    .A2(_14510_),
    .B1(_14511_),
    .Y(_14512_));
 sky130_fd_sc_hd__and3_2 _36871_ (.A(_14506_),
    .B(_14507_),
    .C(_14508_),
    .X(_14513_));
 sky130_fd_sc_hd__nand2_1 _36872_ (.A(_14509_),
    .B(_14511_),
    .Y(_14514_));
 sky130_fd_sc_hd__nor2_2 _36873_ (.A(_14513_),
    .B(_14514_),
    .Y(_14515_));
 sky130_fd_sc_hd__o2bb2ai_4 _36874_ (.A1_N(_14475_),
    .A2_N(_14480_),
    .B1(_14512_),
    .B2(_14515_),
    .Y(_14516_));
 sky130_fd_sc_hd__a21oi_1 _36875_ (.A1(_14506_),
    .A2(_14507_),
    .B1(_14508_),
    .Y(_14517_));
 sky130_fd_sc_hd__o21ai_1 _36876_ (.A1(_14517_),
    .A2(_14513_),
    .B1(_14511_),
    .Y(_14518_));
 sky130_fd_sc_hd__nand3b_1 _36877_ (.A_N(_14511_),
    .B(_14509_),
    .C(_14510_),
    .Y(_14519_));
 sky130_fd_sc_hd__nand2_2 _36878_ (.A(_14518_),
    .B(_14519_),
    .Y(_14520_));
 sky130_fd_sc_hd__nand3_4 _36879_ (.A(_14520_),
    .B(_14480_),
    .C(_14475_),
    .Y(_14521_));
 sky130_vsdinv _36880_ (.A(_14112_),
    .Y(_14522_));
 sky130_fd_sc_hd__o21ai_2 _36881_ (.A1(_14044_),
    .A2(_14047_),
    .B1(_14114_),
    .Y(_14523_));
 sky130_fd_sc_hd__o2bb2ai_4 _36882_ (.A1_N(_14160_),
    .A2_N(_14120_),
    .B1(_14522_),
    .B2(_14523_),
    .Y(_14524_));
 sky130_fd_sc_hd__a21oi_4 _36883_ (.A1(_14516_),
    .A2(_14521_),
    .B1(_14524_),
    .Y(_14525_));
 sky130_fd_sc_hd__and3_1 _36884_ (.A(_14410_),
    .B(_14469_),
    .C(_14474_),
    .X(_14526_));
 sky130_fd_sc_hd__nand2_1 _36885_ (.A(_14520_),
    .B(_14480_),
    .Y(_14527_));
 sky130_fd_sc_hd__o211a_2 _36886_ (.A1(_14526_),
    .A2(_14527_),
    .B1(_14524_),
    .C1(_14516_),
    .X(_14528_));
 sky130_fd_sc_hd__o22ai_4 _36887_ (.A1(_14406_),
    .A2(_14408_),
    .B1(_14525_),
    .B2(_14528_),
    .Y(_14529_));
 sky130_fd_sc_hd__a21oi_2 _36888_ (.A1(_14157_),
    .A2(_14161_),
    .B1(_14043_),
    .Y(_14530_));
 sky130_fd_sc_hd__o21ai_4 _36889_ (.A1(_14247_),
    .A2(_14530_),
    .B1(_14162_),
    .Y(_14531_));
 sky130_fd_sc_hd__a21o_2 _36890_ (.A1(_14516_),
    .A2(_14521_),
    .B1(_14524_),
    .X(_14532_));
 sky130_fd_sc_hd__nand3_4 _36891_ (.A(_14516_),
    .B(_14524_),
    .C(_14521_),
    .Y(_14533_));
 sky130_fd_sc_hd__nor2_8 _36892_ (.A(_14408_),
    .B(_14406_),
    .Y(_14534_));
 sky130_fd_sc_hd__nand3_4 _36893_ (.A(_14532_),
    .B(_14533_),
    .C(_14534_),
    .Y(_14535_));
 sky130_fd_sc_hd__nand3_4 _36894_ (.A(_14529_),
    .B(_14531_),
    .C(_14535_),
    .Y(_14536_));
 sky130_fd_sc_hd__o21ai_2 _36895_ (.A1(_14525_),
    .A2(_14528_),
    .B1(_14534_),
    .Y(_14537_));
 sky130_fd_sc_hd__a21boi_4 _36896_ (.A1(_14242_),
    .A2(_14167_),
    .B1_N(_14162_),
    .Y(_14538_));
 sky130_fd_sc_hd__a21o_1 _36897_ (.A1(_14405_),
    .A2(_14402_),
    .B1(_14407_),
    .X(_14539_));
 sky130_fd_sc_hd__nand3_1 _36898_ (.A(_14405_),
    .B(_14402_),
    .C(_14407_),
    .Y(_14540_));
 sky130_fd_sc_hd__nand2_1 _36899_ (.A(_14539_),
    .B(_14540_),
    .Y(_14541_));
 sky130_fd_sc_hd__nand3_2 _36900_ (.A(_14532_),
    .B(_14533_),
    .C(_14541_),
    .Y(_14542_));
 sky130_fd_sc_hd__nand3_4 _36901_ (.A(_14537_),
    .B(_14538_),
    .C(_14542_),
    .Y(_14543_));
 sky130_fd_sc_hd__a21oi_4 _36902_ (.A1(_14209_),
    .A2(_14210_),
    .B1(_14206_),
    .Y(_14544_));
 sky130_fd_sc_hd__nor2_2 _36903_ (.A(_14211_),
    .B(_14544_),
    .Y(_14545_));
 sky130_fd_sc_hd__nand3_4 _36904_ (.A(_14545_),
    .B(_13944_),
    .C(_13946_),
    .Y(_14546_));
 sky130_fd_sc_hd__o211ai_4 _36905_ (.A1(_14211_),
    .A2(_14544_),
    .B1(_13953_),
    .C1(_13951_),
    .Y(_14547_));
 sky130_fd_sc_hd__buf_2 _36906_ (.A(_14256_),
    .X(_14548_));
 sky130_fd_sc_hd__a21oi_2 _36907_ (.A1(_14546_),
    .A2(_14547_),
    .B1(_14548_),
    .Y(_14549_));
 sky130_fd_sc_hd__and3_1 _36908_ (.A(_14546_),
    .B(_14547_),
    .C(_14256_),
    .X(_14550_));
 sky130_fd_sc_hd__a21oi_2 _36909_ (.A1(_14205_),
    .A2(_14221_),
    .B1(_14204_),
    .Y(_14551_));
 sky130_fd_sc_hd__o21ai_4 _36910_ (.A1(_14549_),
    .A2(_14550_),
    .B1(_14551_),
    .Y(_14552_));
 sky130_fd_sc_hd__o22ai_4 _36911_ (.A1(_14225_),
    .A2(_14226_),
    .B1(_14217_),
    .B2(_14214_),
    .Y(_14553_));
 sky130_fd_sc_hd__nand3_2 _36912_ (.A(_14546_),
    .B(_14547_),
    .C(_14257_),
    .Y(_14554_));
 sky130_fd_sc_hd__a21o_1 _36913_ (.A1(_14546_),
    .A2(_14547_),
    .B1(_14548_),
    .X(_14555_));
 sky130_fd_sc_hd__nand3_4 _36914_ (.A(_14553_),
    .B(_14554_),
    .C(_14555_),
    .Y(_14556_));
 sky130_vsdinv _36915_ (.A(_14256_),
    .Y(_14557_));
 sky130_fd_sc_hd__o21ai_4 _36916_ (.A1(_14557_),
    .A2(_14263_),
    .B1(_14255_),
    .Y(_14558_));
 sky130_fd_sc_hd__a21oi_2 _36917_ (.A1(_14552_),
    .A2(_14556_),
    .B1(_14558_),
    .Y(_14559_));
 sky130_vsdinv _36918_ (.A(_14255_),
    .Y(_14560_));
 sky130_fd_sc_hd__nor2_1 _36919_ (.A(_14557_),
    .B(_14263_),
    .Y(_14561_));
 sky130_fd_sc_hd__o211a_1 _36920_ (.A1(_14560_),
    .A2(_14561_),
    .B1(_14556_),
    .C1(_14552_),
    .X(_14562_));
 sky130_fd_sc_hd__o21a_1 _36921_ (.A1(_14267_),
    .A2(_14262_),
    .B1(_14270_),
    .X(_14563_));
 sky130_fd_sc_hd__o21ai_4 _36922_ (.A1(_14559_),
    .A2(_14562_),
    .B1(_14563_),
    .Y(_14564_));
 sky130_fd_sc_hd__a21o_1 _36923_ (.A1(_14552_),
    .A2(_14556_),
    .B1(_14558_),
    .X(_14565_));
 sky130_fd_sc_hd__o21ai_2 _36924_ (.A1(_14267_),
    .A2(_14262_),
    .B1(_14270_),
    .Y(_14566_));
 sky130_fd_sc_hd__nand3_2 _36925_ (.A(_14552_),
    .B(_14556_),
    .C(_14558_),
    .Y(_14567_));
 sky130_fd_sc_hd__nand3_4 _36926_ (.A(_14565_),
    .B(_14566_),
    .C(_14567_),
    .Y(_14568_));
 sky130_fd_sc_hd__a21oi_2 _36927_ (.A1(_14564_),
    .A2(_14568_),
    .B1(_13663_),
    .Y(_14569_));
 sky130_fd_sc_hd__and3_1 _36928_ (.A(_14564_),
    .B(_13978_),
    .C(_14568_),
    .X(_14570_));
 sky130_fd_sc_hd__nand2_1 _36929_ (.A(_14231_),
    .B(_14234_),
    .Y(_14571_));
 sky130_fd_sc_hd__a21oi_2 _36930_ (.A1(_13879_),
    .A2(_13917_),
    .B1(_14237_),
    .Y(_14572_));
 sky130_fd_sc_hd__a21oi_2 _36931_ (.A1(_14234_),
    .A2(_14235_),
    .B1(_14231_),
    .Y(_14573_));
 sky130_fd_sc_hd__o22ai_4 _36932_ (.A1(_14229_),
    .A2(_14571_),
    .B1(_14572_),
    .B2(_14573_),
    .Y(_14574_));
 sky130_fd_sc_hd__o21bai_4 _36933_ (.A1(_14569_),
    .A2(_14570_),
    .B1_N(_14574_),
    .Y(_14575_));
 sky130_vsdinv _36934_ (.A(_14568_),
    .Y(_14576_));
 sky130_fd_sc_hd__nand2_2 _36935_ (.A(_14564_),
    .B(_13978_),
    .Y(_14577_));
 sky130_fd_sc_hd__a21o_1 _36936_ (.A1(_14564_),
    .A2(_14568_),
    .B1(_13978_),
    .X(_14578_));
 sky130_fd_sc_hd__o211ai_4 _36937_ (.A1(_14576_),
    .A2(_14577_),
    .B1(_14574_),
    .C1(_14578_),
    .Y(_14579_));
 sky130_fd_sc_hd__nor2_1 _36938_ (.A(_13655_),
    .B(_14274_),
    .Y(_14580_));
 sky130_fd_sc_hd__or2_2 _36939_ (.A(_14278_),
    .B(_14580_),
    .X(_14581_));
 sky130_fd_sc_hd__a21oi_4 _36940_ (.A1(_14575_),
    .A2(_14579_),
    .B1(_14581_),
    .Y(_14582_));
 sky130_fd_sc_hd__o211a_1 _36941_ (.A1(_14278_),
    .A2(_14580_),
    .B1(_14579_),
    .C1(_14575_),
    .X(_14583_));
 sky130_fd_sc_hd__o2bb2ai_4 _36942_ (.A1_N(_14536_),
    .A2_N(_14543_),
    .B1(_14582_),
    .B2(_14583_),
    .Y(_14584_));
 sky130_fd_sc_hd__nor2_2 _36943_ (.A(_14582_),
    .B(_14583_),
    .Y(_14585_));
 sky130_fd_sc_hd__nand3_4 _36944_ (.A(_14585_),
    .B(_14536_),
    .C(_14543_),
    .Y(_14586_));
 sky130_vsdinv _36945_ (.A(_14243_),
    .Y(_14587_));
 sky130_fd_sc_hd__nand3_2 _36946_ (.A(_14241_),
    .B(_13931_),
    .C(_14040_),
    .Y(_14588_));
 sky130_fd_sc_hd__o22ai_4 _36947_ (.A1(_14587_),
    .A2(_14588_),
    .B1(_14299_),
    .B2(_14244_),
    .Y(_14589_));
 sky130_fd_sc_hd__a21o_2 _36948_ (.A1(_14584_),
    .A2(_14586_),
    .B1(_14589_),
    .X(_14590_));
 sky130_fd_sc_hd__nand3_4 _36949_ (.A(_14584_),
    .B(_14589_),
    .C(_14586_),
    .Y(_14591_));
 sky130_fd_sc_hd__buf_6 _36950_ (.A(_14305_),
    .X(_14592_));
 sky130_fd_sc_hd__nand2_4 _36951_ (.A(_14298_),
    .B(_14290_),
    .Y(_14593_));
 sky130_fd_sc_hd__nor2_4 _36952_ (.A(_14592_),
    .B(_14593_),
    .Y(_14594_));
 sky130_fd_sc_hd__buf_6 _36953_ (.A(_13719_),
    .X(_14595_));
 sky130_vsdinv _36954_ (.A(_14593_),
    .Y(_14596_));
 sky130_fd_sc_hd__nor2_8 _36955_ (.A(_14595_),
    .B(_14596_),
    .Y(_14597_));
 sky130_fd_sc_hd__nor2_4 _36956_ (.A(_14594_),
    .B(_14597_),
    .Y(_14598_));
 sky130_fd_sc_hd__nand3_4 _36957_ (.A(_14590_),
    .B(_14591_),
    .C(_14598_),
    .Y(_14599_));
 sky130_fd_sc_hd__a21oi_4 _36958_ (.A1(_14584_),
    .A2(_14586_),
    .B1(_14589_),
    .Y(_14600_));
 sky130_fd_sc_hd__and3_1 _36959_ (.A(_14529_),
    .B(_14531_),
    .C(_14535_),
    .X(_14601_));
 sky130_fd_sc_hd__nand2_1 _36960_ (.A(_14575_),
    .B(_14579_),
    .Y(_14602_));
 sky130_fd_sc_hd__nor2_1 _36961_ (.A(_14278_),
    .B(_14580_),
    .Y(_14603_));
 sky130_fd_sc_hd__nand2_1 _36962_ (.A(_14602_),
    .B(_14603_),
    .Y(_14604_));
 sky130_fd_sc_hd__nand3_4 _36963_ (.A(_14581_),
    .B(_14575_),
    .C(_14579_),
    .Y(_14605_));
 sky130_fd_sc_hd__nand3_2 _36964_ (.A(_14543_),
    .B(_14604_),
    .C(_14605_),
    .Y(_14606_));
 sky130_fd_sc_hd__o211a_4 _36965_ (.A1(_14601_),
    .A2(_14606_),
    .B1(_14589_),
    .C1(_14584_),
    .X(_14607_));
 sky130_fd_sc_hd__o22ai_4 _36966_ (.A1(_14597_),
    .A2(_14594_),
    .B1(_14600_),
    .B2(_14607_),
    .Y(_14608_));
 sky130_fd_sc_hd__o211ai_4 _36967_ (.A1(_14324_),
    .A2(_14310_),
    .B1(_14599_),
    .C1(_14608_),
    .Y(_14609_));
 sky130_fd_sc_hd__nor2_4 _36968_ (.A(_14592_),
    .B(_14596_),
    .Y(_14610_));
 sky130_fd_sc_hd__nor2_4 _36969_ (.A(_14595_),
    .B(_14593_),
    .Y(_14611_));
 sky130_fd_sc_hd__o22ai_4 _36970_ (.A1(_14610_),
    .A2(_14611_),
    .B1(_14600_),
    .B2(_14607_),
    .Y(_14612_));
 sky130_fd_sc_hd__a21oi_4 _36971_ (.A1(_14317_),
    .A2(_14322_),
    .B1(_14324_),
    .Y(_14613_));
 sky130_fd_sc_hd__nor2_2 _36972_ (.A(_14611_),
    .B(_14610_),
    .Y(_14614_));
 sky130_fd_sc_hd__nand3_2 _36973_ (.A(_14590_),
    .B(_14591_),
    .C(_14614_),
    .Y(_14615_));
 sky130_fd_sc_hd__nand3_4 _36974_ (.A(_14612_),
    .B(_14613_),
    .C(_14615_),
    .Y(_14616_));
 sky130_fd_sc_hd__a21oi_2 _36975_ (.A1(_14609_),
    .A2(_14616_),
    .B1(_14319_),
    .Y(_14617_));
 sky130_fd_sc_hd__and3_1 _36976_ (.A(_14609_),
    .B(_14616_),
    .C(_14319_),
    .X(_14618_));
 sky130_fd_sc_hd__a21boi_2 _36977_ (.A1(_14328_),
    .A2(_13722_),
    .B1_N(_14321_),
    .Y(_14619_));
 sky130_fd_sc_hd__o21ai_4 _36978_ (.A1(_14617_),
    .A2(_14618_),
    .B1(_14619_),
    .Y(_14620_));
 sky130_vsdinv _36979_ (.A(_13722_),
    .Y(_14621_));
 sky130_fd_sc_hd__a21oi_1 _36980_ (.A1(_14320_),
    .A2(_14316_),
    .B1(_14036_),
    .Y(_14622_));
 sky130_fd_sc_hd__o21ai_2 _36981_ (.A1(_14621_),
    .A2(_14622_),
    .B1(_14321_),
    .Y(_14623_));
 sky130_fd_sc_hd__nand3_2 _36982_ (.A(_14609_),
    .B(_14616_),
    .C(_14319_),
    .Y(_14624_));
 sky130_fd_sc_hd__a21o_1 _36983_ (.A1(_14609_),
    .A2(_14616_),
    .B1(_14319_),
    .X(_14625_));
 sky130_fd_sc_hd__nand3_4 _36984_ (.A(_14623_),
    .B(_14624_),
    .C(_14625_),
    .Y(_14626_));
 sky130_fd_sc_hd__nand2_2 _36985_ (.A(_14620_),
    .B(_14626_),
    .Y(_14627_));
 sky130_fd_sc_hd__nand2_1 _36986_ (.A(_14339_),
    .B(_14024_),
    .Y(_14628_));
 sky130_fd_sc_hd__nand2_1 _36987_ (.A(_14628_),
    .B(_14338_),
    .Y(_14629_));
 sky130_fd_sc_hd__a21bo_2 _36988_ (.A1(_14034_),
    .A2(_14340_),
    .B1_N(_14629_),
    .X(_14630_));
 sky130_fd_sc_hd__xnor2_4 _36989_ (.A(_14627_),
    .B(_14630_),
    .Y(_02661_));
 sky130_fd_sc_hd__a21oi_4 _36990_ (.A1(_14590_),
    .A2(_14598_),
    .B1(_14607_),
    .Y(_14631_));
 sky130_fd_sc_hd__nand2_2 _36991_ (.A(_14605_),
    .B(_14579_),
    .Y(_14632_));
 sky130_vsdinv _36992_ (.A(_14632_),
    .Y(_14633_));
 sky130_fd_sc_hd__nor2_4 _36993_ (.A(_14305_),
    .B(_14633_),
    .Y(_14634_));
 sky130_fd_sc_hd__nor2_4 _36994_ (.A(_14595_),
    .B(_14632_),
    .Y(_14635_));
 sky130_fd_sc_hd__o21ai_2 _36995_ (.A1(_14541_),
    .A2(_14525_),
    .B1(_14533_),
    .Y(_14636_));
 sky130_fd_sc_hd__and3_1 _36996_ (.A(_14436_),
    .B(_14440_),
    .C(_14437_),
    .X(_14637_));
 sky130_fd_sc_hd__a31oi_4 _36997_ (.A1(_14442_),
    .A2(_14446_),
    .A3(_14445_),
    .B1(_14472_),
    .Y(_14638_));
 sky130_fd_sc_hd__nand2_1 _36998_ (.A(_09722_),
    .B(_07343_),
    .Y(_14639_));
 sky130_fd_sc_hd__nand2_4 _36999_ (.A(_10257_),
    .B(_07067_),
    .Y(_14640_));
 sky130_fd_sc_hd__or2_4 _37000_ (.A(_14639_),
    .B(_14640_),
    .X(_14641_));
 sky130_fd_sc_hd__nor2_2 _37001_ (.A(_08578_),
    .B(_10960_),
    .Y(_14642_));
 sky130_fd_sc_hd__nand2_1 _37002_ (.A(_14639_),
    .B(_14640_),
    .Y(_14643_));
 sky130_fd_sc_hd__nand3_4 _37003_ (.A(_14641_),
    .B(_14642_),
    .C(_14643_),
    .Y(_14644_));
 sky130_fd_sc_hd__a31o_2 _37004_ (.A1(_14428_),
    .A2(_19592_),
    .A3(_19885_),
    .B1(_14427_),
    .X(_14645_));
 sky130_fd_sc_hd__a21o_1 _37005_ (.A1(_14084_),
    .A2(_14452_),
    .B1(_14639_),
    .X(_14646_));
 sky130_fd_sc_hd__a21o_1 _37006_ (.A1(_14087_),
    .A2(_07344_),
    .B1(_14640_),
    .X(_14647_));
 sky130_fd_sc_hd__nand3b_4 _37007_ (.A_N(_14642_),
    .B(_14646_),
    .C(_14647_),
    .Y(_14648_));
 sky130_fd_sc_hd__nand3_4 _37008_ (.A(_14644_),
    .B(_14645_),
    .C(_14648_),
    .Y(_14649_));
 sky130_fd_sc_hd__o21a_2 _37009_ (.A1(_14448_),
    .A2(_14450_),
    .B1(_14457_),
    .X(_14650_));
 sky130_fd_sc_hd__a21oi_4 _37010_ (.A1(_14644_),
    .A2(_14648_),
    .B1(_14645_),
    .Y(_14651_));
 sky130_fd_sc_hd__nor2_4 _37011_ (.A(_14650_),
    .B(_14651_),
    .Y(_14652_));
 sky130_fd_sc_hd__nor2_1 _37012_ (.A(_14427_),
    .B(_14430_),
    .Y(_14653_));
 sky130_fd_sc_hd__o2bb2ai_1 _37013_ (.A1_N(_14648_),
    .A2_N(_14644_),
    .B1(_14429_),
    .B2(_14653_),
    .Y(_14654_));
 sky130_fd_sc_hd__a21boi_4 _37014_ (.A1(_14654_),
    .A2(_14649_),
    .B1_N(_14650_),
    .Y(_14655_));
 sky130_fd_sc_hd__a21oi_4 _37015_ (.A1(_14649_),
    .A2(_14652_),
    .B1(_14655_),
    .Y(_14656_));
 sky130_fd_sc_hd__o21a_1 _37016_ (.A1(_14435_),
    .A2(_14422_),
    .B1(_14439_),
    .X(_14657_));
 sky130_fd_sc_hd__nand2_2 _37017_ (.A(_11348_),
    .B(_06464_),
    .Y(_14658_));
 sky130_fd_sc_hd__nand2_2 _37018_ (.A(_10046_),
    .B(_07322_),
    .Y(_14659_));
 sky130_fd_sc_hd__nor2_4 _37019_ (.A(_14658_),
    .B(_14659_),
    .Y(_14660_));
 sky130_fd_sc_hd__and2_1 _37020_ (.A(_14658_),
    .B(_14659_),
    .X(_14661_));
 sky130_fd_sc_hd__nand2_2 _37021_ (.A(_10251_),
    .B(_07052_),
    .Y(_14662_));
 sky130_vsdinv _37022_ (.A(_14662_),
    .Y(_14663_));
 sky130_fd_sc_hd__o21a_1 _37023_ (.A1(_14660_),
    .A2(_14661_),
    .B1(_14663_),
    .X(_14664_));
 sky130_vsdinv _37024_ (.A(_14660_),
    .Y(_14665_));
 sky130_fd_sc_hd__nand2_1 _37025_ (.A(_14658_),
    .B(_14659_),
    .Y(_14666_));
 sky130_fd_sc_hd__and3_1 _37026_ (.A(_14665_),
    .B(_14662_),
    .C(_14666_),
    .X(_14667_));
 sky130_fd_sc_hd__nand3_4 _37027_ (.A(_12780_),
    .B(_19576_),
    .C(_06788_),
    .Y(_14668_));
 sky130_fd_sc_hd__nor2_4 _37028_ (.A(_10365_),
    .B(_14668_),
    .Y(_14669_));
 sky130_fd_sc_hd__nand2_1 _37029_ (.A(_12401_),
    .B(_06650_),
    .Y(_14670_));
 sky130_fd_sc_hd__o21a_1 _37030_ (.A1(_10365_),
    .A2(_18474_),
    .B1(_14670_),
    .X(_14671_));
 sky130_fd_sc_hd__o22ai_4 _37031_ (.A1(_10286_),
    .A2(_07275_),
    .B1(_14669_),
    .B2(_14671_),
    .Y(_14672_));
 sky130_fd_sc_hd__nor2_4 _37032_ (.A(_10286_),
    .B(_07275_),
    .Y(_14673_));
 sky130_fd_sc_hd__o21ai_2 _37033_ (.A1(_10365_),
    .A2(_13745_),
    .B1(_14670_),
    .Y(_14674_));
 sky130_fd_sc_hd__nand3b_4 _37034_ (.A_N(_14669_),
    .B(_14673_),
    .C(_14674_),
    .Y(_14675_));
 sky130_fd_sc_hd__o21ai_4 _37035_ (.A1(_14414_),
    .A2(_14413_),
    .B1(_14417_),
    .Y(_14676_));
 sky130_fd_sc_hd__a21oi_4 _37036_ (.A1(_14672_),
    .A2(_14675_),
    .B1(_14676_),
    .Y(_14677_));
 sky130_fd_sc_hd__o21ai_1 _37037_ (.A1(_19899_),
    .A2(_14668_),
    .B1(_14673_),
    .Y(_14678_));
 sky130_fd_sc_hd__o211a_2 _37038_ (.A1(_14671_),
    .A2(_14678_),
    .B1(_14676_),
    .C1(_14672_),
    .X(_14679_));
 sky130_fd_sc_hd__o22ai_4 _37039_ (.A1(_14664_),
    .A2(_14667_),
    .B1(_14677_),
    .B2(_14679_),
    .Y(_14680_));
 sky130_fd_sc_hd__a21o_1 _37040_ (.A1(_14672_),
    .A2(_14675_),
    .B1(_14676_),
    .X(_14681_));
 sky130_fd_sc_hd__nand3_4 _37041_ (.A(_14672_),
    .B(_14675_),
    .C(_14676_),
    .Y(_14682_));
 sky130_fd_sc_hd__nand3_2 _37042_ (.A(_14665_),
    .B(_14663_),
    .C(_14666_),
    .Y(_14683_));
 sky130_fd_sc_hd__o21ai_1 _37043_ (.A1(_14660_),
    .A2(_14661_),
    .B1(_14662_),
    .Y(_14684_));
 sky130_fd_sc_hd__nand2_2 _37044_ (.A(_14683_),
    .B(_14684_),
    .Y(_14685_));
 sky130_fd_sc_hd__nand3_2 _37045_ (.A(_14681_),
    .B(_14682_),
    .C(_14685_),
    .Y(_14686_));
 sky130_fd_sc_hd__nand3_4 _37046_ (.A(_14657_),
    .B(_14680_),
    .C(_14686_),
    .Y(_14687_));
 sky130_vsdinv _37047_ (.A(_14684_),
    .Y(_14688_));
 sky130_vsdinv _37048_ (.A(_14683_),
    .Y(_14689_));
 sky130_fd_sc_hd__o22ai_4 _37049_ (.A1(_14688_),
    .A2(_14689_),
    .B1(_14677_),
    .B2(_14679_),
    .Y(_14690_));
 sky130_fd_sc_hd__nand3b_2 _37050_ (.A_N(_14685_),
    .B(_14681_),
    .C(_14682_),
    .Y(_14691_));
 sky130_fd_sc_hd__o21ai_2 _37051_ (.A1(_14435_),
    .A2(_14422_),
    .B1(_14439_),
    .Y(_14692_));
 sky130_fd_sc_hd__nand3_4 _37052_ (.A(_14690_),
    .B(_14691_),
    .C(_14692_),
    .Y(_14693_));
 sky130_fd_sc_hd__nand3_2 _37053_ (.A(_14656_),
    .B(_14687_),
    .C(_14693_),
    .Y(_14694_));
 sky130_fd_sc_hd__and2_1 _37054_ (.A(_14652_),
    .B(_14649_),
    .X(_14695_));
 sky130_fd_sc_hd__o2bb2ai_1 _37055_ (.A1_N(_14693_),
    .A2_N(_14687_),
    .B1(_14655_),
    .B2(_14695_),
    .Y(_14696_));
 sky130_fd_sc_hd__o211ai_4 _37056_ (.A1(_14637_),
    .A2(_14638_),
    .B1(_14694_),
    .C1(_14696_),
    .Y(_14697_));
 sky130_fd_sc_hd__nand2_1 _37057_ (.A(_14687_),
    .B(_14693_),
    .Y(_14698_));
 sky130_fd_sc_hd__nand2_4 _37058_ (.A(_14698_),
    .B(_14656_),
    .Y(_14699_));
 sky130_fd_sc_hd__nand2_1 _37059_ (.A(_14441_),
    .B(_14472_),
    .Y(_14700_));
 sky130_fd_sc_hd__nand2_2 _37060_ (.A(_14700_),
    .B(_14447_),
    .Y(_14701_));
 sky130_fd_sc_hd__a21o_1 _37061_ (.A1(_14649_),
    .A2(_14652_),
    .B1(_14655_),
    .X(_14702_));
 sky130_fd_sc_hd__nand3_4 _37062_ (.A(_14702_),
    .B(_14687_),
    .C(_14693_),
    .Y(_14703_));
 sky130_fd_sc_hd__nand3_4 _37063_ (.A(_14699_),
    .B(_14701_),
    .C(_14703_),
    .Y(_14704_));
 sky130_fd_sc_hd__nor2_2 _37064_ (.A(_14463_),
    .B(_14466_),
    .Y(_14705_));
 sky130_fd_sc_hd__a21oi_4 _37065_ (.A1(_14489_),
    .A2(_14488_),
    .B1(_14483_),
    .Y(_14706_));
 sky130_fd_sc_hd__nand2_4 _37066_ (.A(_08908_),
    .B(_07701_),
    .Y(_14707_));
 sky130_fd_sc_hd__nand2_4 _37067_ (.A(_08541_),
    .B(_08333_),
    .Y(_14708_));
 sky130_fd_sc_hd__nor2_8 _37068_ (.A(_14707_),
    .B(_14708_),
    .Y(_14709_));
 sky130_fd_sc_hd__and2_1 _37069_ (.A(_14707_),
    .B(_14708_),
    .X(_14710_));
 sky130_fd_sc_hd__nand2_2 _37070_ (.A(_12470_),
    .B(_10458_),
    .Y(_14711_));
 sky130_fd_sc_hd__o21ai_2 _37071_ (.A1(_14709_),
    .A2(_14710_),
    .B1(_14711_),
    .Y(_14712_));
 sky130_vsdinv _37072_ (.A(_14711_),
    .Y(_14713_));
 sky130_fd_sc_hd__nand2_4 _37073_ (.A(_14707_),
    .B(_14708_),
    .Y(_14714_));
 sky130_fd_sc_hd__nand3b_4 _37074_ (.A_N(_14709_),
    .B(_14713_),
    .C(_14714_),
    .Y(_14715_));
 sky130_fd_sc_hd__nand3b_4 _37075_ (.A_N(_14706_),
    .B(_14712_),
    .C(_14715_),
    .Y(_14716_));
 sky130_fd_sc_hd__o21ai_2 _37076_ (.A1(_14709_),
    .A2(_14710_),
    .B1(_14713_),
    .Y(_14717_));
 sky130_fd_sc_hd__nand3b_2 _37077_ (.A_N(_14709_),
    .B(_14711_),
    .C(_14714_),
    .Y(_14718_));
 sky130_fd_sc_hd__nand3_4 _37078_ (.A(_14717_),
    .B(_14718_),
    .C(_14706_),
    .Y(_14719_));
 sky130_fd_sc_hd__nand2_2 _37079_ (.A(_07484_),
    .B(_10459_),
    .Y(_14720_));
 sky130_fd_sc_hd__nand2_4 _37080_ (.A(_07825_),
    .B(_19854_),
    .Y(_14721_));
 sky130_fd_sc_hd__nor2_4 _37081_ (.A(_14720_),
    .B(_14721_),
    .Y(_14722_));
 sky130_fd_sc_hd__and2_1 _37082_ (.A(_14720_),
    .B(_14721_),
    .X(_14723_));
 sky130_fd_sc_hd__nor2_1 _37083_ (.A(_14722_),
    .B(_14723_),
    .Y(_14724_));
 sky130_fd_sc_hd__nor2_4 _37084_ (.A(net471),
    .B(_11537_),
    .Y(_14725_));
 sky130_vsdinv _37085_ (.A(_14725_),
    .Y(_14726_));
 sky130_fd_sc_hd__nand2_1 _37086_ (.A(_14724_),
    .B(_14726_),
    .Y(_14727_));
 sky130_fd_sc_hd__o21ai_1 _37087_ (.A1(_14722_),
    .A2(_14723_),
    .B1(_14725_),
    .Y(_14728_));
 sky130_fd_sc_hd__nand2_2 _37088_ (.A(_14727_),
    .B(_14728_),
    .Y(_14729_));
 sky130_fd_sc_hd__a21oi_2 _37089_ (.A1(_14716_),
    .A2(_14719_),
    .B1(_14729_),
    .Y(_14730_));
 sky130_fd_sc_hd__nor3_2 _37090_ (.A(_14722_),
    .B(_14725_),
    .C(_14723_),
    .Y(_14731_));
 sky130_fd_sc_hd__nor2_1 _37091_ (.A(_14726_),
    .B(_14724_),
    .Y(_14732_));
 sky130_fd_sc_hd__o211a_1 _37092_ (.A1(_14731_),
    .A2(_14732_),
    .B1(_14716_),
    .C1(_14719_),
    .X(_14733_));
 sky130_fd_sc_hd__o22ai_4 _37093_ (.A1(_14470_),
    .A2(_14705_),
    .B1(_14730_),
    .B2(_14733_),
    .Y(_14734_));
 sky130_fd_sc_hd__nand2_4 _37094_ (.A(_14467_),
    .B(_14462_),
    .Y(_14735_));
 sky130_fd_sc_hd__a21o_1 _37095_ (.A1(_14716_),
    .A2(_14719_),
    .B1(_14729_),
    .X(_14736_));
 sky130_fd_sc_hd__nand3_4 _37096_ (.A(_14729_),
    .B(_14716_),
    .C(_14719_),
    .Y(_14737_));
 sky130_fd_sc_hd__nand3_4 _37097_ (.A(_14735_),
    .B(_14736_),
    .C(_14737_),
    .Y(_14738_));
 sky130_fd_sc_hd__nand2_1 _37098_ (.A(_14505_),
    .B(_14495_),
    .Y(_14739_));
 sky130_fd_sc_hd__nand2_1 _37099_ (.A(_14739_),
    .B(_14491_),
    .Y(_14740_));
 sky130_vsdinv _37100_ (.A(_14740_),
    .Y(_14741_));
 sky130_fd_sc_hd__nand3_2 _37101_ (.A(_14734_),
    .B(_14738_),
    .C(_14741_),
    .Y(_14742_));
 sky130_vsdinv _37102_ (.A(_14742_),
    .Y(_14743_));
 sky130_fd_sc_hd__a21o_1 _37103_ (.A1(_14734_),
    .A2(_14738_),
    .B1(_14741_),
    .X(_14744_));
 sky130_vsdinv _37104_ (.A(_14744_),
    .Y(_14745_));
 sky130_fd_sc_hd__o2bb2ai_1 _37105_ (.A1_N(_14697_),
    .A2_N(_14704_),
    .B1(_14743_),
    .B2(_14745_),
    .Y(_14746_));
 sky130_fd_sc_hd__a21boi_4 _37106_ (.A1(_14520_),
    .A2(_14480_),
    .B1_N(_14475_),
    .Y(_14747_));
 sky130_vsdinv _37107_ (.A(_14495_),
    .Y(_14748_));
 sky130_fd_sc_hd__and3_1 _37108_ (.A(_14491_),
    .B(_14503_),
    .C(_14504_),
    .X(_14749_));
 sky130_fd_sc_hd__o2bb2ai_1 _37109_ (.A1_N(_14738_),
    .A2_N(_14734_),
    .B1(_14748_),
    .B2(_14749_),
    .Y(_14750_));
 sky130_fd_sc_hd__nand3_1 _37110_ (.A(_14734_),
    .B(_14738_),
    .C(_14740_),
    .Y(_14751_));
 sky130_fd_sc_hd__nand2_1 _37111_ (.A(_14750_),
    .B(_14751_),
    .Y(_14752_));
 sky130_fd_sc_hd__nand3_2 _37112_ (.A(_14704_),
    .B(_14697_),
    .C(_14752_),
    .Y(_14753_));
 sky130_fd_sc_hd__nand3_4 _37113_ (.A(_14746_),
    .B(_14747_),
    .C(_14753_),
    .Y(_14754_));
 sky130_fd_sc_hd__nand2_2 _37114_ (.A(_14527_),
    .B(_14475_),
    .Y(_14755_));
 sky130_vsdinv _37115_ (.A(_14751_),
    .Y(_14756_));
 sky130_vsdinv _37116_ (.A(_14750_),
    .Y(_14757_));
 sky130_fd_sc_hd__o2bb2ai_2 _37117_ (.A1_N(_14697_),
    .A2_N(_14704_),
    .B1(_14756_),
    .B2(_14757_),
    .Y(_14758_));
 sky130_fd_sc_hd__nand2_2 _37118_ (.A(_14744_),
    .B(_14742_),
    .Y(_14759_));
 sky130_fd_sc_hd__nand3_4 _37119_ (.A(_14759_),
    .B(_14704_),
    .C(_14697_),
    .Y(_14760_));
 sky130_fd_sc_hd__nand3_4 _37120_ (.A(_14755_),
    .B(_14758_),
    .C(_14760_),
    .Y(_14761_));
 sky130_fd_sc_hd__o21a_2 _37121_ (.A1(_14395_),
    .A2(_14367_),
    .B1(_14400_),
    .X(_14762_));
 sky130_fd_sc_hd__nand2_1 _37122_ (.A(_14514_),
    .B(_14510_),
    .Y(_14763_));
 sky130_fd_sc_hd__nand2_1 _37123_ (.A(_08615_),
    .B(_19848_),
    .Y(_14764_));
 sky130_fd_sc_hd__nand2_1 _37124_ (.A(_08616_),
    .B(_09950_),
    .Y(_14765_));
 sky130_fd_sc_hd__or2_2 _37125_ (.A(_14764_),
    .B(_14765_),
    .X(_14766_));
 sky130_fd_sc_hd__nor2_2 _37126_ (.A(net444),
    .B(_09805_),
    .Y(_14767_));
 sky130_fd_sc_hd__nand2_1 _37127_ (.A(_14764_),
    .B(_14765_),
    .Y(_14768_));
 sky130_fd_sc_hd__nand3_4 _37128_ (.A(_14766_),
    .B(_14767_),
    .C(_14768_),
    .Y(_14769_));
 sky130_fd_sc_hd__a21o_1 _37129_ (.A1(_19637_),
    .A2(_10493_),
    .B1(_14764_),
    .X(_14770_));
 sky130_fd_sc_hd__a21o_1 _37130_ (.A1(_19633_),
    .A2(_19849_),
    .B1(_14765_),
    .X(_14771_));
 sky130_fd_sc_hd__nand3b_4 _37131_ (.A_N(_14767_),
    .B(_14770_),
    .C(_14771_),
    .Y(_14772_));
 sky130_fd_sc_hd__a31o_2 _37132_ (.A1(_14499_),
    .A2(_13408_),
    .A3(_19856_),
    .B1(_14498_),
    .X(_14773_));
 sky130_fd_sc_hd__a21oi_4 _37133_ (.A1(_14769_),
    .A2(_14772_),
    .B1(_14773_),
    .Y(_14774_));
 sky130_fd_sc_hd__a21oi_1 _37134_ (.A1(_14496_),
    .A2(_14497_),
    .B1(_14502_),
    .Y(_14775_));
 sky130_fd_sc_hd__o211a_1 _37135_ (.A1(_14498_),
    .A2(_14775_),
    .B1(_14772_),
    .C1(_14769_),
    .X(_14776_));
 sky130_fd_sc_hd__nand2_2 _37136_ (.A(_14353_),
    .B(_14350_),
    .Y(_14777_));
 sky130_vsdinv _37137_ (.A(_14777_),
    .Y(_14778_));
 sky130_fd_sc_hd__o21ai_4 _37138_ (.A1(_14774_),
    .A2(_14776_),
    .B1(_14778_),
    .Y(_14779_));
 sky130_fd_sc_hd__a21o_1 _37139_ (.A1(_14769_),
    .A2(_14772_),
    .B1(_14773_),
    .X(_14780_));
 sky130_fd_sc_hd__nand3_4 _37140_ (.A(_14769_),
    .B(_14773_),
    .C(_14772_),
    .Y(_14781_));
 sky130_fd_sc_hd__nand3_4 _37141_ (.A(_14780_),
    .B(_14781_),
    .C(_14777_),
    .Y(_14782_));
 sky130_fd_sc_hd__o21ai_4 _37142_ (.A1(_14364_),
    .A2(_14357_),
    .B1(_14363_),
    .Y(_14783_));
 sky130_fd_sc_hd__a21oi_4 _37143_ (.A1(_14779_),
    .A2(_14782_),
    .B1(_14783_),
    .Y(_14784_));
 sky130_fd_sc_hd__and3_1 _37144_ (.A(_14779_),
    .B(_14782_),
    .C(_14783_),
    .X(_14785_));
 sky130_fd_sc_hd__nor2_2 _37145_ (.A(_14371_),
    .B(_14373_),
    .Y(_14786_));
 sky130_fd_sc_hd__a21oi_4 _37146_ (.A1(_14377_),
    .A2(_14378_),
    .B1(_14786_),
    .Y(_14787_));
 sky130_fd_sc_hd__nor2_2 _37147_ (.A(_11721_),
    .B(_12618_),
    .Y(_14788_));
 sky130_fd_sc_hd__nand2_2 _37148_ (.A(_06896_),
    .B(_09933_),
    .Y(_14789_));
 sky130_fd_sc_hd__a21o_1 _37149_ (.A1(_06343_),
    .A2(_11199_),
    .B1(_14789_),
    .X(_14790_));
 sky130_fd_sc_hd__nand2_2 _37150_ (.A(_19647_),
    .B(_19829_),
    .Y(_14791_));
 sky130_fd_sc_hd__a21o_1 _37151_ (.A1(_06342_),
    .A2(_10598_),
    .B1(_14791_),
    .X(_14792_));
 sky130_fd_sc_hd__nand3b_4 _37152_ (.A_N(_14788_),
    .B(_14790_),
    .C(_14792_),
    .Y(_14793_));
 sky130_fd_sc_hd__nand3_2 _37153_ (.A(_08597_),
    .B(_09439_),
    .C(_10487_),
    .Y(_14794_));
 sky130_fd_sc_hd__nand2_1 _37154_ (.A(_14789_),
    .B(_14791_),
    .Y(_14795_));
 sky130_fd_sc_hd__o211ai_4 _37155_ (.A1(_10597_),
    .A2(_14794_),
    .B1(_14795_),
    .C1(_14788_),
    .Y(_14796_));
 sky130_fd_sc_hd__nand2_2 _37156_ (.A(_14793_),
    .B(_14796_),
    .Y(_14797_));
 sky130_fd_sc_hd__nor2_4 _37157_ (.A(_14787_),
    .B(_14797_),
    .Y(_14798_));
 sky130_fd_sc_hd__nand2_2 _37158_ (.A(_14797_),
    .B(_14787_),
    .Y(_14799_));
 sky130_vsdinv _37159_ (.A(_06018_),
    .Y(_14800_));
 sky130_fd_sc_hd__o21a_2 _37160_ (.A1(_06401_),
    .A2(_05882_),
    .B1(_11184_),
    .X(_14801_));
 sky130_fd_sc_hd__o21ai_4 _37161_ (.A1(_14800_),
    .A2(_14385_),
    .B1(_14801_),
    .Y(_14802_));
 sky130_fd_sc_hd__nor2_4 _37162_ (.A(_05616_),
    .B(_14802_),
    .Y(_14803_));
 sky130_fd_sc_hd__o21ai_2 _37163_ (.A1(_06018_),
    .A2(_05736_),
    .B1(_11593_),
    .Y(_14804_));
 sky130_fd_sc_hd__and3_4 _37164_ (.A(_12274_),
    .B(_19651_),
    .C(_06158_),
    .X(_14805_));
 sky130_fd_sc_hd__nor2_2 _37165_ (.A(_14804_),
    .B(_14805_),
    .Y(_14806_));
 sky130_fd_sc_hd__nor2_4 _37166_ (.A(_14207_),
    .B(_14806_),
    .Y(_14807_));
 sky130_fd_sc_hd__nor2_2 _37167_ (.A(_14803_),
    .B(_14807_),
    .Y(_14808_));
 sky130_fd_sc_hd__buf_4 _37168_ (.A(_14808_),
    .X(_14809_));
 sky130_fd_sc_hd__nand3b_2 _37169_ (.A_N(_14798_),
    .B(_14799_),
    .C(_14809_),
    .Y(_14810_));
 sky130_fd_sc_hd__a31o_1 _37170_ (.A1(_14378_),
    .A2(net478),
    .A3(_19830_),
    .B1(_14786_),
    .X(_14811_));
 sky130_fd_sc_hd__a21oi_4 _37171_ (.A1(_14793_),
    .A2(_14796_),
    .B1(_14811_),
    .Y(_14812_));
 sky130_fd_sc_hd__nand2_1 _37172_ (.A(_14802_),
    .B(_14206_),
    .Y(_14813_));
 sky130_fd_sc_hd__o21ai_2 _37173_ (.A1(_05616_),
    .A2(_14802_),
    .B1(_14813_),
    .Y(_14814_));
 sky130_fd_sc_hd__buf_6 _37174_ (.A(_14814_),
    .X(_14815_));
 sky130_fd_sc_hd__o21ai_2 _37175_ (.A1(_14812_),
    .A2(_14798_),
    .B1(_14815_),
    .Y(_14816_));
 sky130_fd_sc_hd__nand2_4 _37176_ (.A(_14810_),
    .B(_14816_),
    .Y(_14817_));
 sky130_fd_sc_hd__o21ai_2 _37177_ (.A1(_14784_),
    .A2(_14785_),
    .B1(_14817_),
    .Y(_14818_));
 sky130_fd_sc_hd__a21o_1 _37178_ (.A1(_14779_),
    .A2(_14782_),
    .B1(_14783_),
    .X(_14819_));
 sky130_fd_sc_hd__nand3_4 _37179_ (.A(_14779_),
    .B(_14782_),
    .C(_14783_),
    .Y(_14820_));
 sky130_fd_sc_hd__nand3b_2 _37180_ (.A_N(_14817_),
    .B(_14819_),
    .C(_14820_),
    .Y(_14821_));
 sky130_fd_sc_hd__nand3_4 _37181_ (.A(_14763_),
    .B(_14818_),
    .C(_14821_),
    .Y(_14822_));
 sky130_fd_sc_hd__o21bai_4 _37182_ (.A1(_14784_),
    .A2(_14785_),
    .B1_N(_14817_),
    .Y(_14823_));
 sky130_fd_sc_hd__a21oi_4 _37183_ (.A1(_14509_),
    .A2(_14511_),
    .B1(_14513_),
    .Y(_14824_));
 sky130_fd_sc_hd__nand3_4 _37184_ (.A(_14819_),
    .B(_14817_),
    .C(_14820_),
    .Y(_14825_));
 sky130_fd_sc_hd__nand3_4 _37185_ (.A(_14823_),
    .B(_14824_),
    .C(_14825_),
    .Y(_14826_));
 sky130_fd_sc_hd__nand2_1 _37186_ (.A(_14822_),
    .B(_14826_),
    .Y(_14827_));
 sky130_fd_sc_hd__nor2_1 _37187_ (.A(_14762_),
    .B(_14827_),
    .Y(_14828_));
 sky130_vsdinv _37188_ (.A(_14762_),
    .Y(_14829_));
 sky130_fd_sc_hd__a21oi_4 _37189_ (.A1(_14822_),
    .A2(_14826_),
    .B1(_14829_),
    .Y(_14830_));
 sky130_fd_sc_hd__o2bb2ai_2 _37190_ (.A1_N(_14754_),
    .A2_N(_14761_),
    .B1(_14828_),
    .B2(_14830_),
    .Y(_14831_));
 sky130_fd_sc_hd__a31oi_4 _37191_ (.A1(_14823_),
    .A2(_14824_),
    .A3(_14825_),
    .B1(_14762_),
    .Y(_14832_));
 sky130_fd_sc_hd__a21oi_4 _37192_ (.A1(_14822_),
    .A2(_14832_),
    .B1(_14830_),
    .Y(_14833_));
 sky130_fd_sc_hd__nand3_4 _37193_ (.A(_14833_),
    .B(_14754_),
    .C(_14761_),
    .Y(_14834_));
 sky130_fd_sc_hd__nand3_4 _37194_ (.A(_14636_),
    .B(_14831_),
    .C(_14834_),
    .Y(_14835_));
 sky130_fd_sc_hd__a21oi_4 _37195_ (.A1(_14532_),
    .A2(_14534_),
    .B1(_14528_),
    .Y(_14836_));
 sky130_fd_sc_hd__nand2_1 _37196_ (.A(_14827_),
    .B(_14762_),
    .Y(_14837_));
 sky130_fd_sc_hd__nand2_1 _37197_ (.A(_14832_),
    .B(_14822_),
    .Y(_14838_));
 sky130_fd_sc_hd__nand2_1 _37198_ (.A(_14837_),
    .B(_14838_),
    .Y(_14839_));
 sky130_fd_sc_hd__nand3_2 _37199_ (.A(_14839_),
    .B(_14754_),
    .C(_14761_),
    .Y(_14840_));
 sky130_fd_sc_hd__nand2_1 _37200_ (.A(_14761_),
    .B(_14754_),
    .Y(_14841_));
 sky130_fd_sc_hd__nand2_1 _37201_ (.A(_14841_),
    .B(_14833_),
    .Y(_14842_));
 sky130_fd_sc_hd__nand3_4 _37202_ (.A(_14836_),
    .B(_14840_),
    .C(_14842_),
    .Y(_14843_));
 sky130_fd_sc_hd__a21oi_4 _37203_ (.A1(_14384_),
    .A2(_14385_),
    .B1(_14206_),
    .Y(_14844_));
 sky130_fd_sc_hd__nor2_2 _37204_ (.A(_14386_),
    .B(_14844_),
    .Y(_14845_));
 sky130_fd_sc_hd__nand3_4 _37205_ (.A(_14845_),
    .B(_13944_),
    .C(_13946_),
    .Y(_14846_));
 sky130_fd_sc_hd__o211ai_4 _37206_ (.A1(_14386_),
    .A2(_14844_),
    .B1(_13953_),
    .C1(_13951_),
    .Y(_14847_));
 sky130_fd_sc_hd__a21o_1 _37207_ (.A1(_14846_),
    .A2(_14847_),
    .B1(_14548_),
    .X(_14848_));
 sky130_fd_sc_hd__nand3_4 _37208_ (.A(_14846_),
    .B(_14847_),
    .C(_14548_),
    .Y(_14849_));
 sky130_fd_sc_hd__nand2_2 _37209_ (.A(_14848_),
    .B(_14849_),
    .Y(_14850_));
 sky130_fd_sc_hd__nor2_4 _37210_ (.A(_14381_),
    .B(_14380_),
    .Y(_14851_));
 sky130_fd_sc_hd__nor2_4 _37211_ (.A(_14851_),
    .B(_14393_),
    .Y(_14852_));
 sky130_fd_sc_hd__nand2_4 _37212_ (.A(_14850_),
    .B(_14852_),
    .Y(_14853_));
 sky130_fd_sc_hd__o211ai_4 _37213_ (.A1(_14851_),
    .A2(_14393_),
    .B1(_14849_),
    .C1(_14848_),
    .Y(_14854_));
 sky130_fd_sc_hd__nand2_1 _37214_ (.A(_14853_),
    .B(_14854_),
    .Y(_14855_));
 sky130_vsdinv _37215_ (.A(_14547_),
    .Y(_14856_));
 sky130_fd_sc_hd__a21oi_2 _37216_ (.A1(_14548_),
    .A2(_14546_),
    .B1(_14856_),
    .Y(_14857_));
 sky130_fd_sc_hd__nand2_2 _37217_ (.A(_14855_),
    .B(_14857_),
    .Y(_14858_));
 sky130_vsdinv _37218_ (.A(_14857_),
    .Y(_14859_));
 sky130_fd_sc_hd__nand3_4 _37219_ (.A(_14853_),
    .B(_14854_),
    .C(_14859_),
    .Y(_14860_));
 sky130_fd_sc_hd__nand2_1 _37220_ (.A(_14552_),
    .B(_14558_),
    .Y(_14861_));
 sky130_fd_sc_hd__nand2_4 _37221_ (.A(_14861_),
    .B(_14556_),
    .Y(_14862_));
 sky130_fd_sc_hd__a21oi_4 _37222_ (.A1(_14858_),
    .A2(_14860_),
    .B1(_14862_),
    .Y(_14863_));
 sky130_fd_sc_hd__and3_1 _37223_ (.A(_14858_),
    .B(_14862_),
    .C(_14860_),
    .X(_14864_));
 sky130_fd_sc_hd__o21ai_2 _37224_ (.A1(_14863_),
    .A2(_14864_),
    .B1(_13663_),
    .Y(_14865_));
 sky130_fd_sc_hd__a21oi_2 _37225_ (.A1(_14396_),
    .A2(_14401_),
    .B1(_14397_),
    .Y(_14866_));
 sky130_fd_sc_hd__a21oi_4 _37226_ (.A1(_14402_),
    .A2(_14407_),
    .B1(_14866_),
    .Y(_14867_));
 sky130_fd_sc_hd__a21oi_1 _37227_ (.A1(_14853_),
    .A2(_14854_),
    .B1(_14859_),
    .Y(_14868_));
 sky130_fd_sc_hd__and3_1 _37228_ (.A(_14853_),
    .B(_14854_),
    .C(_14859_),
    .X(_14869_));
 sky130_fd_sc_hd__o21bai_2 _37229_ (.A1(_14868_),
    .A2(_14869_),
    .B1_N(_14862_),
    .Y(_14870_));
 sky130_fd_sc_hd__nand3_4 _37230_ (.A(_14858_),
    .B(_14862_),
    .C(_14860_),
    .Y(_14871_));
 sky130_fd_sc_hd__nand3_2 _37231_ (.A(_14870_),
    .B(_13655_),
    .C(_14871_),
    .Y(_14872_));
 sky130_fd_sc_hd__nand3_4 _37232_ (.A(_14865_),
    .B(_14867_),
    .C(_14872_),
    .Y(_14873_));
 sky130_fd_sc_hd__o2bb2ai_1 _37233_ (.A1_N(_14871_),
    .A2_N(_14870_),
    .B1(_13653_),
    .B2(_13651_),
    .Y(_14874_));
 sky130_fd_sc_hd__nand2_1 _37234_ (.A(_14402_),
    .B(_14407_),
    .Y(_14875_));
 sky130_fd_sc_hd__nand2_1 _37235_ (.A(_14875_),
    .B(_14405_),
    .Y(_14876_));
 sky130_fd_sc_hd__nand3_2 _37236_ (.A(_14870_),
    .B(_13978_),
    .C(_14871_),
    .Y(_14877_));
 sky130_fd_sc_hd__nand3_4 _37237_ (.A(_14874_),
    .B(_14876_),
    .C(_14877_),
    .Y(_14878_));
 sky130_fd_sc_hd__nand2_2 _37238_ (.A(_14577_),
    .B(_14568_),
    .Y(_14879_));
 sky130_fd_sc_hd__a21oi_4 _37239_ (.A1(_14873_),
    .A2(_14878_),
    .B1(_14879_),
    .Y(_14880_));
 sky130_vsdinv _37240_ (.A(_14564_),
    .Y(_14881_));
 sky130_fd_sc_hd__nor2_1 _37241_ (.A(_14283_),
    .B(_14881_),
    .Y(_14882_));
 sky130_fd_sc_hd__o211a_2 _37242_ (.A1(_14576_),
    .A2(_14882_),
    .B1(_14878_),
    .C1(_14873_),
    .X(_14883_));
 sky130_fd_sc_hd__o2bb2ai_4 _37243_ (.A1_N(_14835_),
    .A2_N(_14843_),
    .B1(_14880_),
    .B2(_14883_),
    .Y(_14884_));
 sky130_fd_sc_hd__nor2_4 _37244_ (.A(_14880_),
    .B(_14883_),
    .Y(_14885_));
 sky130_fd_sc_hd__nand3_4 _37245_ (.A(_14885_),
    .B(_14843_),
    .C(_14835_),
    .Y(_14886_));
 sky130_vsdinv _37246_ (.A(_14535_),
    .Y(_14887_));
 sky130_fd_sc_hd__nand2_1 _37247_ (.A(_14529_),
    .B(_14531_),
    .Y(_14888_));
 sky130_fd_sc_hd__nand2_1 _37248_ (.A(_14604_),
    .B(_14605_),
    .Y(_14889_));
 sky130_fd_sc_hd__a21oi_2 _37249_ (.A1(_14529_),
    .A2(_14535_),
    .B1(_14531_),
    .Y(_14890_));
 sky130_fd_sc_hd__o22ai_4 _37250_ (.A1(_14887_),
    .A2(_14888_),
    .B1(_14889_),
    .B2(_14890_),
    .Y(_14891_));
 sky130_fd_sc_hd__a21oi_4 _37251_ (.A1(_14884_),
    .A2(_14886_),
    .B1(_14891_),
    .Y(_14892_));
 sky130_vsdinv _37252_ (.A(_14835_),
    .Y(_14893_));
 sky130_fd_sc_hd__nand2_2 _37253_ (.A(_14885_),
    .B(_14843_),
    .Y(_14894_));
 sky130_fd_sc_hd__o211a_2 _37254_ (.A1(_14893_),
    .A2(_14894_),
    .B1(_14884_),
    .C1(_14891_),
    .X(_14895_));
 sky130_fd_sc_hd__o22ai_4 _37255_ (.A1(_14634_),
    .A2(_14635_),
    .B1(_14892_),
    .B2(_14895_),
    .Y(_14896_));
 sky130_fd_sc_hd__a21o_1 _37256_ (.A1(_14884_),
    .A2(_14886_),
    .B1(_14891_),
    .X(_14897_));
 sky130_fd_sc_hd__nand3_4 _37257_ (.A(_14891_),
    .B(_14884_),
    .C(_14886_),
    .Y(_14898_));
 sky130_fd_sc_hd__nor2_4 _37258_ (.A(_14635_),
    .B(_14634_),
    .Y(_14899_));
 sky130_fd_sc_hd__nand3_2 _37259_ (.A(_14897_),
    .B(_14898_),
    .C(_14899_),
    .Y(_14900_));
 sky130_fd_sc_hd__nand3_4 _37260_ (.A(_14631_),
    .B(_14896_),
    .C(_14900_),
    .Y(_14901_));
 sky130_fd_sc_hd__nor2_8 _37261_ (.A(_14329_),
    .B(_14633_),
    .Y(_14902_));
 sky130_fd_sc_hd__buf_6 _37262_ (.A(_14592_),
    .X(_14903_));
 sky130_fd_sc_hd__nor2_2 _37263_ (.A(_14903_),
    .B(_14632_),
    .Y(_14904_));
 sky130_fd_sc_hd__o22ai_4 _37264_ (.A1(_14902_),
    .A2(_14904_),
    .B1(_14892_),
    .B2(_14895_),
    .Y(_14905_));
 sky130_fd_sc_hd__o21ai_2 _37265_ (.A1(_14614_),
    .A2(_14600_),
    .B1(_14591_),
    .Y(_14906_));
 sky130_fd_sc_hd__nand3b_4 _37266_ (.A_N(_14899_),
    .B(_14897_),
    .C(_14898_),
    .Y(_14907_));
 sky130_fd_sc_hd__nand3_4 _37267_ (.A(_14905_),
    .B(_14906_),
    .C(_14907_),
    .Y(_14908_));
 sky130_fd_sc_hd__nand3_4 _37268_ (.A(_14901_),
    .B(_14908_),
    .C(_14597_),
    .Y(_14909_));
 sky130_vsdinv _37269_ (.A(_14909_),
    .Y(_14910_));
 sky130_fd_sc_hd__o2bb2ai_4 _37270_ (.A1_N(_14908_),
    .A2_N(_14901_),
    .B1(_14331_),
    .B2(_14596_),
    .Y(_14911_));
 sky130_fd_sc_hd__nand2_1 _37271_ (.A(_14616_),
    .B(_14319_),
    .Y(_14912_));
 sky130_fd_sc_hd__nand2_1 _37272_ (.A(_14912_),
    .B(_14609_),
    .Y(_14913_));
 sky130_fd_sc_hd__nand2_2 _37273_ (.A(_14911_),
    .B(_14913_),
    .Y(_14914_));
 sky130_fd_sc_hd__a21o_1 _37274_ (.A1(_14911_),
    .A2(_14909_),
    .B1(_14913_),
    .X(_14915_));
 sky130_fd_sc_hd__o21a_2 _37275_ (.A1(_14910_),
    .A2(_14914_),
    .B1(_14915_),
    .X(_14916_));
 sky130_fd_sc_hd__a21bo_1 _37276_ (.A1(_14630_),
    .A2(_14620_),
    .B1_N(_14626_),
    .X(_14917_));
 sky130_fd_sc_hd__xor2_4 _37277_ (.A(_14916_),
    .B(_14917_),
    .X(_02662_));
 sky130_fd_sc_hd__nand2_2 _37278_ (.A(_06924_),
    .B(_19843_),
    .Y(_14918_));
 sky130_fd_sc_hd__nand2_2 _37279_ (.A(_08623_),
    .B(_10488_),
    .Y(_14919_));
 sky130_fd_sc_hd__nor2_2 _37280_ (.A(_14918_),
    .B(_14919_),
    .Y(_14920_));
 sky130_fd_sc_hd__and2_1 _37281_ (.A(_14918_),
    .B(_14919_),
    .X(_14921_));
 sky130_fd_sc_hd__nor2_2 _37282_ (.A(net444),
    .B(_11206_),
    .Y(_14922_));
 sky130_fd_sc_hd__o21bai_4 _37283_ (.A1(_14920_),
    .A2(_14921_),
    .B1_N(_14922_),
    .Y(_14923_));
 sky130_fd_sc_hd__or2_2 _37284_ (.A(_14918_),
    .B(_14919_),
    .X(_14924_));
 sky130_fd_sc_hd__nand2_1 _37285_ (.A(_14918_),
    .B(_14919_),
    .Y(_14925_));
 sky130_fd_sc_hd__nand3_4 _37286_ (.A(_14924_),
    .B(_14922_),
    .C(_14925_),
    .Y(_14926_));
 sky130_fd_sc_hd__nand2_2 _37287_ (.A(_14720_),
    .B(_14721_),
    .Y(_14927_));
 sky130_fd_sc_hd__a31o_2 _37288_ (.A1(_14927_),
    .A2(_19629_),
    .A3(_19853_),
    .B1(_14722_),
    .X(_14928_));
 sky130_fd_sc_hd__a21oi_4 _37289_ (.A1(_14923_),
    .A2(_14926_),
    .B1(_14928_),
    .Y(_14929_));
 sky130_fd_sc_hd__a21oi_4 _37290_ (.A1(_14725_),
    .A2(_14927_),
    .B1(_14722_),
    .Y(_14930_));
 sky130_fd_sc_hd__nand2_2 _37291_ (.A(_14923_),
    .B(_14926_),
    .Y(_14931_));
 sky130_fd_sc_hd__nor2_4 _37292_ (.A(_14930_),
    .B(_14931_),
    .Y(_14932_));
 sky130_fd_sc_hd__and2_2 _37293_ (.A(_14769_),
    .B(_14766_),
    .X(_14933_));
 sky130_fd_sc_hd__o21ai_4 _37294_ (.A1(_14929_),
    .A2(_14932_),
    .B1(_14933_),
    .Y(_14934_));
 sky130_fd_sc_hd__nand2_2 _37295_ (.A(_14931_),
    .B(_14930_),
    .Y(_14935_));
 sky130_fd_sc_hd__nand3_4 _37296_ (.A(_14923_),
    .B(_14926_),
    .C(_14928_),
    .Y(_14936_));
 sky130_fd_sc_hd__nand2_2 _37297_ (.A(_14769_),
    .B(_14766_),
    .Y(_14937_));
 sky130_fd_sc_hd__nand3_4 _37298_ (.A(_14935_),
    .B(_14936_),
    .C(_14937_),
    .Y(_14938_));
 sky130_fd_sc_hd__o21ai_4 _37299_ (.A1(_14774_),
    .A2(_14778_),
    .B1(_14781_),
    .Y(_14939_));
 sky130_fd_sc_hd__a21oi_4 _37300_ (.A1(_14934_),
    .A2(_14938_),
    .B1(_14939_),
    .Y(_14940_));
 sky130_fd_sc_hd__nand2_1 _37301_ (.A(_14935_),
    .B(_14937_),
    .Y(_14941_));
 sky130_fd_sc_hd__o211a_2 _37302_ (.A1(_14932_),
    .A2(_14941_),
    .B1(_14939_),
    .C1(_14934_),
    .X(_14942_));
 sky130_fd_sc_hd__nand2_2 _37303_ (.A(_08597_),
    .B(_11202_),
    .Y(_14943_));
 sky130_fd_sc_hd__nand2_2 _37304_ (.A(_09439_),
    .B(_19825_),
    .Y(_14944_));
 sky130_fd_sc_hd__nor2_2 _37305_ (.A(_14943_),
    .B(_14944_),
    .Y(_14945_));
 sky130_fd_sc_hd__nand2_2 _37306_ (.A(_12614_),
    .B(_06349_),
    .Y(_14946_));
 sky130_vsdinv _37307_ (.A(_14946_),
    .Y(_14947_));
 sky130_fd_sc_hd__nand2_2 _37308_ (.A(_14943_),
    .B(_14944_),
    .Y(_14948_));
 sky130_fd_sc_hd__nand3b_4 _37309_ (.A_N(_14945_),
    .B(_14947_),
    .C(_14948_),
    .Y(_14949_));
 sky130_fd_sc_hd__a21o_1 _37310_ (.A1(_19648_),
    .A2(_11200_),
    .B1(_14943_),
    .X(_14950_));
 sky130_fd_sc_hd__a21o_1 _37311_ (.A1(_19645_),
    .A2(_19830_),
    .B1(_14944_),
    .X(_14951_));
 sky130_fd_sc_hd__nand3_4 _37312_ (.A(_14950_),
    .B(_14951_),
    .C(_14946_),
    .Y(_14952_));
 sky130_fd_sc_hd__o21ai_4 _37313_ (.A1(_14789_),
    .A2(_14791_),
    .B1(_14796_),
    .Y(_14953_));
 sky130_fd_sc_hd__a21o_2 _37314_ (.A1(_14949_),
    .A2(_14952_),
    .B1(_14953_),
    .X(_14954_));
 sky130_fd_sc_hd__nand3_4 _37315_ (.A(_14953_),
    .B(_14952_),
    .C(_14949_),
    .Y(_14955_));
 sky130_fd_sc_hd__a21oi_4 _37316_ (.A1(_14954_),
    .A2(_14955_),
    .B1(_14809_),
    .Y(_14956_));
 sky130_fd_sc_hd__nand3_4 _37317_ (.A(_14954_),
    .B(_14808_),
    .C(_14955_),
    .Y(_14957_));
 sky130_vsdinv _37318_ (.A(_14957_),
    .Y(_14958_));
 sky130_fd_sc_hd__nor2_4 _37319_ (.A(_14956_),
    .B(_14958_),
    .Y(_14959_));
 sky130_fd_sc_hd__o21ai_4 _37320_ (.A1(_14940_),
    .A2(_14942_),
    .B1(_14959_),
    .Y(_14960_));
 sky130_fd_sc_hd__a21oi_4 _37321_ (.A1(_14736_),
    .A2(_14737_),
    .B1(_14735_),
    .Y(_14961_));
 sky130_fd_sc_hd__o21a_2 _37322_ (.A1(_14741_),
    .A2(_14961_),
    .B1(_14738_),
    .X(_14962_));
 sky130_fd_sc_hd__a21o_1 _37323_ (.A1(_14934_),
    .A2(_14938_),
    .B1(_14939_),
    .X(_14963_));
 sky130_fd_sc_hd__nand3_4 _37324_ (.A(_14934_),
    .B(_14939_),
    .C(_14938_),
    .Y(_14964_));
 sky130_fd_sc_hd__or2b_4 _37325_ (.A(_14956_),
    .B_N(_14957_),
    .X(_14965_));
 sky130_fd_sc_hd__nand3_4 _37326_ (.A(_14963_),
    .B(_14964_),
    .C(_14965_),
    .Y(_14966_));
 sky130_fd_sc_hd__nand3_4 _37327_ (.A(_14960_),
    .B(_14962_),
    .C(_14966_),
    .Y(_14967_));
 sky130_fd_sc_hd__o22ai_4 _37328_ (.A1(_14956_),
    .A2(_14958_),
    .B1(_14940_),
    .B2(_14942_),
    .Y(_14968_));
 sky130_fd_sc_hd__nand3_2 _37329_ (.A(_14963_),
    .B(_14964_),
    .C(_14959_),
    .Y(_14969_));
 sky130_fd_sc_hd__o21ai_2 _37330_ (.A1(_14741_),
    .A2(_14961_),
    .B1(_14738_),
    .Y(_14970_));
 sky130_fd_sc_hd__nand3_4 _37331_ (.A(_14968_),
    .B(_14969_),
    .C(_14970_),
    .Y(_14971_));
 sky130_fd_sc_hd__o21a_1 _37332_ (.A1(_14817_),
    .A2(_14784_),
    .B1(_14820_),
    .X(_14972_));
 sky130_vsdinv _37333_ (.A(_14972_),
    .Y(_14973_));
 sky130_fd_sc_hd__and3_1 _37334_ (.A(_14967_),
    .B(_14971_),
    .C(_14973_),
    .X(_14974_));
 sky130_fd_sc_hd__a21oi_4 _37335_ (.A1(_14967_),
    .A2(_14971_),
    .B1(_14973_),
    .Y(_14975_));
 sky130_fd_sc_hd__nand3_4 _37336_ (.A(_12780_),
    .B(_19576_),
    .C(_06462_),
    .Y(_14976_));
 sky130_fd_sc_hd__nor2_4 _37337_ (.A(_19895_),
    .B(_14976_),
    .Y(_14977_));
 sky130_fd_sc_hd__o22a_2 _37338_ (.A1(_06289_),
    .A2(_13099_),
    .B1(_11338_),
    .B2(net440),
    .X(_14978_));
 sky130_fd_sc_hd__o22ai_4 _37339_ (.A1(_10286_),
    .A2(_06810_),
    .B1(_14977_),
    .B2(_14978_),
    .Y(_14979_));
 sky130_fd_sc_hd__a22o_2 _37340_ (.A1(_13737_),
    .A2(_06286_),
    .B1(net443),
    .B2(_11292_),
    .X(_14980_));
 sky130_fd_sc_hd__nand2_1 _37341_ (.A(_10828_),
    .B(_07327_),
    .Y(_14981_));
 sky130_vsdinv _37342_ (.A(_14981_),
    .Y(_14982_));
 sky130_fd_sc_hd__nand3b_4 _37343_ (.A_N(_14977_),
    .B(_14980_),
    .C(_14982_),
    .Y(_14983_));
 sky130_fd_sc_hd__a21o_2 _37344_ (.A1(_14674_),
    .A2(_14673_),
    .B1(_14669_),
    .X(_14984_));
 sky130_fd_sc_hd__a21oi_4 _37345_ (.A1(_14979_),
    .A2(_14983_),
    .B1(_14984_),
    .Y(_14985_));
 sky130_fd_sc_hd__o21ai_1 _37346_ (.A1(_19895_),
    .A2(_14976_),
    .B1(_14982_),
    .Y(_14986_));
 sky130_fd_sc_hd__o211a_2 _37347_ (.A1(_14978_),
    .A2(_14986_),
    .B1(_14984_),
    .C1(_14979_),
    .X(_14987_));
 sky130_fd_sc_hd__nand2_2 _37348_ (.A(_10251_),
    .B(_07051_),
    .Y(_14988_));
 sky130_vsdinv _37349_ (.A(_14988_),
    .Y(_14989_));
 sky130_fd_sc_hd__nand2_4 _37350_ (.A(_10281_),
    .B(_19884_),
    .Y(_14990_));
 sky130_fd_sc_hd__nand2_2 _37351_ (.A(_19587_),
    .B(_08280_),
    .Y(_14991_));
 sky130_fd_sc_hd__nor2_4 _37352_ (.A(_14990_),
    .B(_14991_),
    .Y(_14992_));
 sky130_fd_sc_hd__and2_2 _37353_ (.A(_14990_),
    .B(_14991_),
    .X(_14993_));
 sky130_fd_sc_hd__nor3_4 _37354_ (.A(_14989_),
    .B(_14992_),
    .C(_14993_),
    .Y(_14994_));
 sky130_fd_sc_hd__o21a_2 _37355_ (.A1(_14992_),
    .A2(_14993_),
    .B1(_14989_),
    .X(_14995_));
 sky130_fd_sc_hd__nor2_8 _37356_ (.A(_14994_),
    .B(_14995_),
    .Y(_14996_));
 sky130_fd_sc_hd__o21ai_2 _37357_ (.A1(_14985_),
    .A2(_14987_),
    .B1(_14996_),
    .Y(_14997_));
 sky130_fd_sc_hd__o21ai_2 _37358_ (.A1(_14685_),
    .A2(_14677_),
    .B1(_14682_),
    .Y(_14998_));
 sky130_fd_sc_hd__a21o_1 _37359_ (.A1(_14979_),
    .A2(_14983_),
    .B1(_14984_),
    .X(_14999_));
 sky130_fd_sc_hd__nand3_4 _37360_ (.A(_14979_),
    .B(_14984_),
    .C(_14983_),
    .Y(_15000_));
 sky130_fd_sc_hd__nand3b_2 _37361_ (.A_N(_14996_),
    .B(_14999_),
    .C(_15000_),
    .Y(_15001_));
 sky130_fd_sc_hd__nand3_4 _37362_ (.A(_14997_),
    .B(_14998_),
    .C(_15001_),
    .Y(_15002_));
 sky130_fd_sc_hd__o21bai_4 _37363_ (.A1(_14985_),
    .A2(_14987_),
    .B1_N(_14996_),
    .Y(_15003_));
 sky130_fd_sc_hd__o21a_2 _37364_ (.A1(_14685_),
    .A2(_14677_),
    .B1(_14682_),
    .X(_15004_));
 sky130_fd_sc_hd__nand3_4 _37365_ (.A(_14999_),
    .B(_15000_),
    .C(_14996_),
    .Y(_15005_));
 sky130_fd_sc_hd__nand3_4 _37366_ (.A(_15003_),
    .B(_15004_),
    .C(_15005_),
    .Y(_15006_));
 sky130_fd_sc_hd__nand2_1 _37367_ (.A(_10260_),
    .B(_09607_),
    .Y(_15007_));
 sky130_fd_sc_hd__nand2_1 _37368_ (.A(_09723_),
    .B(_07325_),
    .Y(_15008_));
 sky130_fd_sc_hd__or2_2 _37369_ (.A(_15007_),
    .B(_15008_),
    .X(_15009_));
 sky130_fd_sc_hd__nor2_2 _37370_ (.A(_08579_),
    .B(_10654_),
    .Y(_15010_));
 sky130_fd_sc_hd__nand2_1 _37371_ (.A(_15007_),
    .B(_15008_),
    .Y(_15011_));
 sky130_fd_sc_hd__nand3_4 _37372_ (.A(_15009_),
    .B(_15010_),
    .C(_15011_),
    .Y(_15012_));
 sky130_fd_sc_hd__a21o_1 _37373_ (.A1(_14084_),
    .A2(_10957_),
    .B1(_15007_),
    .X(_15013_));
 sky130_fd_sc_hd__a21o_1 _37374_ (.A1(_14087_),
    .A2(_19874_),
    .B1(_15008_),
    .X(_15014_));
 sky130_fd_sc_hd__nand3b_4 _37375_ (.A_N(_15010_),
    .B(_15013_),
    .C(_15014_),
    .Y(_15015_));
 sky130_fd_sc_hd__nand2_2 _37376_ (.A(_15012_),
    .B(_15015_),
    .Y(_15016_));
 sky130_fd_sc_hd__a21o_2 _37377_ (.A1(_14663_),
    .A2(_14666_),
    .B1(_14660_),
    .X(_15017_));
 sky130_vsdinv _37378_ (.A(_15017_),
    .Y(_15018_));
 sky130_fd_sc_hd__nand2_2 _37379_ (.A(_15016_),
    .B(_15018_),
    .Y(_15019_));
 sky130_fd_sc_hd__nand3_4 _37380_ (.A(_15012_),
    .B(_15015_),
    .C(_15017_),
    .Y(_15020_));
 sky130_fd_sc_hd__nand2_2 _37381_ (.A(_14644_),
    .B(_14641_),
    .Y(_15021_));
 sky130_fd_sc_hd__a21oi_4 _37382_ (.A1(_15019_),
    .A2(_15020_),
    .B1(_15021_),
    .Y(_15022_));
 sky130_fd_sc_hd__a21oi_1 _37383_ (.A1(_14658_),
    .A2(_14659_),
    .B1(_14662_),
    .Y(_15023_));
 sky130_fd_sc_hd__o211a_2 _37384_ (.A1(_14660_),
    .A2(_15023_),
    .B1(_15015_),
    .C1(_15012_),
    .X(_15024_));
 sky130_fd_sc_hd__nand2_2 _37385_ (.A(_15019_),
    .B(_15021_),
    .Y(_15025_));
 sky130_fd_sc_hd__nor2_1 _37386_ (.A(_15024_),
    .B(_15025_),
    .Y(_15026_));
 sky130_fd_sc_hd__o2bb2ai_1 _37387_ (.A1_N(_15002_),
    .A2_N(_15006_),
    .B1(_15022_),
    .B2(_15026_),
    .Y(_15027_));
 sky130_fd_sc_hd__nand2_1 _37388_ (.A(_14656_),
    .B(_14687_),
    .Y(_15028_));
 sky130_fd_sc_hd__nand2_1 _37389_ (.A(_15028_),
    .B(_14693_),
    .Y(_15029_));
 sky130_fd_sc_hd__a22oi_4 _37390_ (.A1(_14641_),
    .A2(_14644_),
    .B1(_15016_),
    .B2(_15018_),
    .Y(_15030_));
 sky130_fd_sc_hd__a21oi_4 _37391_ (.A1(_15020_),
    .A2(_15030_),
    .B1(_15022_),
    .Y(_15031_));
 sky130_fd_sc_hd__nand3_2 _37392_ (.A(_15006_),
    .B(_15031_),
    .C(_15002_),
    .Y(_15032_));
 sky130_fd_sc_hd__nand3_4 _37393_ (.A(_15027_),
    .B(_15029_),
    .C(_15032_),
    .Y(_15033_));
 sky130_fd_sc_hd__nand2_1 _37394_ (.A(_15006_),
    .B(_15002_),
    .Y(_15034_));
 sky130_fd_sc_hd__nand2_2 _37395_ (.A(_15034_),
    .B(_15031_),
    .Y(_15035_));
 sky130_fd_sc_hd__a21oi_4 _37396_ (.A1(_15012_),
    .A2(_15015_),
    .B1(_15017_),
    .Y(_15036_));
 sky130_fd_sc_hd__and2_1 _37397_ (.A(_14644_),
    .B(_14641_),
    .X(_15037_));
 sky130_fd_sc_hd__o21ai_2 _37398_ (.A1(_15036_),
    .A2(_15024_),
    .B1(_15037_),
    .Y(_15038_));
 sky130_fd_sc_hd__o21ai_4 _37399_ (.A1(_15024_),
    .A2(_15025_),
    .B1(_15038_),
    .Y(_15039_));
 sky130_fd_sc_hd__nand3_4 _37400_ (.A(_15006_),
    .B(_15002_),
    .C(_15039_),
    .Y(_15040_));
 sky130_fd_sc_hd__a21boi_4 _37401_ (.A1(_14656_),
    .A2(_14687_),
    .B1_N(_14693_),
    .Y(_15041_));
 sky130_fd_sc_hd__nand3_4 _37402_ (.A(_15035_),
    .B(_15040_),
    .C(_15041_),
    .Y(_15042_));
 sky130_fd_sc_hd__nand2_2 _37403_ (.A(_08153_),
    .B(_08333_),
    .Y(_15043_));
 sky130_fd_sc_hd__nand2_2 _37404_ (.A(_08541_),
    .B(_08337_),
    .Y(_15044_));
 sky130_fd_sc_hd__nor2_4 _37405_ (.A(_15043_),
    .B(_15044_),
    .Y(_15045_));
 sky130_fd_sc_hd__and2_1 _37406_ (.A(_15043_),
    .B(_15044_),
    .X(_15046_));
 sky130_fd_sc_hd__nand2_2 _37407_ (.A(_12470_),
    .B(_10459_),
    .Y(_15047_));
 sky130_fd_sc_hd__o21ai_2 _37408_ (.A1(_15045_),
    .A2(_15046_),
    .B1(_15047_),
    .Y(_15048_));
 sky130_fd_sc_hd__nand2_2 _37409_ (.A(_15043_),
    .B(_15044_),
    .Y(_15049_));
 sky130_vsdinv _37410_ (.A(_15047_),
    .Y(_15050_));
 sky130_fd_sc_hd__nand3b_2 _37411_ (.A_N(_15045_),
    .B(_15049_),
    .C(_15050_),
    .Y(_15051_));
 sky130_fd_sc_hd__a21o_1 _37412_ (.A1(_14713_),
    .A2(_14714_),
    .B1(_14709_),
    .X(_15052_));
 sky130_fd_sc_hd__nand3_4 _37413_ (.A(_15048_),
    .B(_15051_),
    .C(_15052_),
    .Y(_15053_));
 sky130_fd_sc_hd__o21ai_2 _37414_ (.A1(_15045_),
    .A2(_15046_),
    .B1(_15050_),
    .Y(_15054_));
 sky130_fd_sc_hd__nand3b_2 _37415_ (.A_N(_15045_),
    .B(_15049_),
    .C(_15047_),
    .Y(_15055_));
 sky130_fd_sc_hd__a21oi_2 _37416_ (.A1(_14713_),
    .A2(_14714_),
    .B1(_14709_),
    .Y(_15056_));
 sky130_fd_sc_hd__nand3_4 _37417_ (.A(_15054_),
    .B(_15055_),
    .C(_15056_),
    .Y(_15057_));
 sky130_fd_sc_hd__nand2_1 _37418_ (.A(_15053_),
    .B(_15057_),
    .Y(_15058_));
 sky130_fd_sc_hd__nand2_2 _37419_ (.A(_07484_),
    .B(_10643_),
    .Y(_15059_));
 sky130_fd_sc_hd__nand2_1 _37420_ (.A(_08565_),
    .B(_19851_),
    .Y(_15060_));
 sky130_fd_sc_hd__nor2_2 _37421_ (.A(_15059_),
    .B(_15060_),
    .Y(_15061_));
 sky130_fd_sc_hd__nand2_1 _37422_ (.A(_15059_),
    .B(_15060_),
    .Y(_15062_));
 sky130_vsdinv _37423_ (.A(_15062_),
    .Y(_15063_));
 sky130_fd_sc_hd__nand2_1 _37424_ (.A(_11003_),
    .B(_19849_),
    .Y(_15064_));
 sky130_fd_sc_hd__o21bai_1 _37425_ (.A1(_15061_),
    .A2(_15063_),
    .B1_N(_15064_),
    .Y(_15065_));
 sky130_fd_sc_hd__nand3b_2 _37426_ (.A_N(_15061_),
    .B(_15064_),
    .C(_15062_),
    .Y(_15066_));
 sky130_fd_sc_hd__and2_1 _37427_ (.A(_15065_),
    .B(_15066_),
    .X(_15067_));
 sky130_fd_sc_hd__nand2_4 _37428_ (.A(_15058_),
    .B(_15067_),
    .Y(_15068_));
 sky130_fd_sc_hd__nand2_2 _37429_ (.A(_15065_),
    .B(_15066_),
    .Y(_15069_));
 sky130_fd_sc_hd__nand3_4 _37430_ (.A(_15069_),
    .B(_15053_),
    .C(_15057_),
    .Y(_15070_));
 sky130_fd_sc_hd__o21ai_4 _37431_ (.A1(_14650_),
    .A2(_14651_),
    .B1(_14649_),
    .Y(_15071_));
 sky130_fd_sc_hd__a21o_1 _37432_ (.A1(_15068_),
    .A2(_15070_),
    .B1(_15071_),
    .X(_15072_));
 sky130_fd_sc_hd__nand3_4 _37433_ (.A(_15071_),
    .B(_15068_),
    .C(_15070_),
    .Y(_15073_));
 sky130_fd_sc_hd__a21bo_1 _37434_ (.A1(_14719_),
    .A2(_14729_),
    .B1_N(_14716_),
    .X(_15074_));
 sky130_fd_sc_hd__a21oi_4 _37435_ (.A1(_15072_),
    .A2(_15073_),
    .B1(_15074_),
    .Y(_15075_));
 sky130_fd_sc_hd__nand3_1 _37436_ (.A(_15072_),
    .B(_15073_),
    .C(_15074_),
    .Y(_15076_));
 sky130_vsdinv _37437_ (.A(_15076_),
    .Y(_15077_));
 sky130_fd_sc_hd__o2bb2ai_4 _37438_ (.A1_N(_15033_),
    .A2_N(_15042_),
    .B1(_15075_),
    .B2(_15077_),
    .Y(_15078_));
 sky130_fd_sc_hd__a21oi_4 _37439_ (.A1(_15068_),
    .A2(_15070_),
    .B1(_15071_),
    .Y(_15079_));
 sky130_vsdinv _37440_ (.A(_15074_),
    .Y(_15080_));
 sky130_fd_sc_hd__nor2_4 _37441_ (.A(_15079_),
    .B(_15080_),
    .Y(_15081_));
 sky130_fd_sc_hd__a21oi_4 _37442_ (.A1(_15073_),
    .A2(_15081_),
    .B1(_15075_),
    .Y(_15082_));
 sky130_fd_sc_hd__nand3_4 _37443_ (.A(_15082_),
    .B(_15042_),
    .C(_15033_),
    .Y(_15083_));
 sky130_fd_sc_hd__a21oi_2 _37444_ (.A1(_14699_),
    .A2(_14703_),
    .B1(_14701_),
    .Y(_15084_));
 sky130_fd_sc_hd__a21o_2 _37445_ (.A1(_14704_),
    .A2(_14759_),
    .B1(_15084_),
    .X(_15085_));
 sky130_fd_sc_hd__a21oi_4 _37446_ (.A1(_15078_),
    .A2(_15083_),
    .B1(_15085_),
    .Y(_15086_));
 sky130_fd_sc_hd__a31oi_1 _37447_ (.A1(_14701_),
    .A2(_14703_),
    .A3(_14699_),
    .B1(_14752_),
    .Y(_15087_));
 sky130_fd_sc_hd__o211a_1 _37448_ (.A1(_15084_),
    .A2(_15087_),
    .B1(_15083_),
    .C1(_15078_),
    .X(_15088_));
 sky130_fd_sc_hd__o22ai_4 _37449_ (.A1(_14974_),
    .A2(_14975_),
    .B1(_15086_),
    .B2(_15088_),
    .Y(_15089_));
 sky130_fd_sc_hd__a21o_1 _37450_ (.A1(_15078_),
    .A2(_15083_),
    .B1(_15085_),
    .X(_15090_));
 sky130_fd_sc_hd__nor2_2 _37451_ (.A(_14975_),
    .B(_14974_),
    .Y(_15091_));
 sky130_fd_sc_hd__nand3_4 _37452_ (.A(_15085_),
    .B(_15078_),
    .C(_15083_),
    .Y(_15092_));
 sky130_fd_sc_hd__nand3_4 _37453_ (.A(_15090_),
    .B(_15091_),
    .C(_15092_),
    .Y(_15093_));
 sky130_fd_sc_hd__a21oi_2 _37454_ (.A1(_14758_),
    .A2(_14760_),
    .B1(_14755_),
    .Y(_15094_));
 sky130_fd_sc_hd__o21ai_2 _37455_ (.A1(_15094_),
    .A2(_14839_),
    .B1(_14761_),
    .Y(_15095_));
 sky130_fd_sc_hd__nand3_4 _37456_ (.A(_15089_),
    .B(_15093_),
    .C(_15095_),
    .Y(_15096_));
 sky130_fd_sc_hd__a21oi_4 _37457_ (.A1(_14960_),
    .A2(_14966_),
    .B1(_14962_),
    .Y(_15097_));
 sky130_fd_sc_hd__nand2_1 _37458_ (.A(_14967_),
    .B(_14973_),
    .Y(_15098_));
 sky130_fd_sc_hd__and2_1 _37459_ (.A(_14817_),
    .B(_14820_),
    .X(_15099_));
 sky130_fd_sc_hd__o2bb2ai_1 _37460_ (.A1_N(_14971_),
    .A2_N(_14967_),
    .B1(_14784_),
    .B2(_15099_),
    .Y(_15100_));
 sky130_fd_sc_hd__o21ai_4 _37461_ (.A1(_15097_),
    .A2(_15098_),
    .B1(_15100_),
    .Y(_15101_));
 sky130_fd_sc_hd__o21bai_2 _37462_ (.A1(_15086_),
    .A2(_15088_),
    .B1_N(_15101_),
    .Y(_15102_));
 sky130_fd_sc_hd__a21boi_4 _37463_ (.A1(_14833_),
    .A2(_14754_),
    .B1_N(_14761_),
    .Y(_15103_));
 sky130_fd_sc_hd__nand3_2 _37464_ (.A(_15090_),
    .B(_15092_),
    .C(_15101_),
    .Y(_15104_));
 sky130_fd_sc_hd__nand3_4 _37465_ (.A(_15102_),
    .B(_15103_),
    .C(_15104_),
    .Y(_15105_));
 sky130_fd_sc_hd__a21oi_4 _37466_ (.A1(_14823_),
    .A2(_14825_),
    .B1(_14824_),
    .Y(_15106_));
 sky130_fd_sc_hd__a21oi_2 _37467_ (.A1(_14826_),
    .A2(_14829_),
    .B1(_15106_),
    .Y(_15107_));
 sky130_fd_sc_hd__nor2_2 _37468_ (.A(_05615_),
    .B(_14804_),
    .Y(_15108_));
 sky130_fd_sc_hd__o211ai_4 _37469_ (.A1(_14805_),
    .A2(_15108_),
    .B1(_13953_),
    .C1(_13951_),
    .Y(_15109_));
 sky130_fd_sc_hd__a21oi_4 _37470_ (.A1(_14801_),
    .A2(_06014_),
    .B1(_14805_),
    .Y(_15110_));
 sky130_fd_sc_hd__nand3_4 _37471_ (.A(_13944_),
    .B(_15110_),
    .C(_13946_),
    .Y(_15111_));
 sky130_fd_sc_hd__nand2_2 _37472_ (.A(_15109_),
    .B(_15111_),
    .Y(_15112_));
 sky130_fd_sc_hd__nand2_8 _37473_ (.A(_15112_),
    .B(_14557_),
    .Y(_15113_));
 sky130_fd_sc_hd__nand3_4 _37474_ (.A(_15109_),
    .B(_15111_),
    .C(_14256_),
    .Y(_15114_));
 sky130_fd_sc_hd__nand2_8 _37475_ (.A(_15113_),
    .B(_15114_),
    .Y(_15115_));
 sky130_fd_sc_hd__a21oi_4 _37476_ (.A1(_14799_),
    .A2(_14809_),
    .B1(_14798_),
    .Y(_15116_));
 sky130_fd_sc_hd__nand2_2 _37477_ (.A(_15115_),
    .B(_15116_),
    .Y(_15117_));
 sky130_vsdinv _37478_ (.A(_14796_),
    .Y(_15118_));
 sky130_fd_sc_hd__nand2_1 _37479_ (.A(_14811_),
    .B(_14793_),
    .Y(_15119_));
 sky130_fd_sc_hd__o22ai_4 _37480_ (.A1(_15118_),
    .A2(_15119_),
    .B1(_14815_),
    .B2(_14812_),
    .Y(_15120_));
 sky130_fd_sc_hd__nand3_4 _37481_ (.A(_15120_),
    .B(_15114_),
    .C(_15113_),
    .Y(_15121_));
 sky130_vsdinv _37482_ (.A(_14847_),
    .Y(_15122_));
 sky130_fd_sc_hd__and2_1 _37483_ (.A(_14846_),
    .B(_14548_),
    .X(_15123_));
 sky130_fd_sc_hd__or2_2 _37484_ (.A(_15122_),
    .B(_15123_),
    .X(_15124_));
 sky130_fd_sc_hd__a21oi_2 _37485_ (.A1(_15117_),
    .A2(_15121_),
    .B1(_15124_),
    .Y(_15125_));
 sky130_fd_sc_hd__o211a_1 _37486_ (.A1(_15122_),
    .A2(_15123_),
    .B1(_15121_),
    .C1(_15117_),
    .X(_15126_));
 sky130_fd_sc_hd__nor2_2 _37487_ (.A(_14852_),
    .B(_14850_),
    .Y(_15127_));
 sky130_fd_sc_hd__a21oi_2 _37488_ (.A1(_14853_),
    .A2(_14859_),
    .B1(_15127_),
    .Y(_15128_));
 sky130_fd_sc_hd__o21ai_4 _37489_ (.A1(_15125_),
    .A2(_15126_),
    .B1(_15128_),
    .Y(_15129_));
 sky130_fd_sc_hd__a21o_1 _37490_ (.A1(_14853_),
    .A2(_14859_),
    .B1(_15127_),
    .X(_15130_));
 sky130_fd_sc_hd__a21o_1 _37491_ (.A1(_15117_),
    .A2(_15121_),
    .B1(_15124_),
    .X(_15131_));
 sky130_fd_sc_hd__nand3_2 _37492_ (.A(_15124_),
    .B(_15117_),
    .C(_15121_),
    .Y(_15132_));
 sky130_fd_sc_hd__nand3_4 _37493_ (.A(_15130_),
    .B(_15131_),
    .C(_15132_),
    .Y(_15133_));
 sky130_fd_sc_hd__a21o_1 _37494_ (.A1(_15129_),
    .A2(_15133_),
    .B1(_13655_),
    .X(_15134_));
 sky130_fd_sc_hd__nand3_2 _37495_ (.A(_15129_),
    .B(_15133_),
    .C(_13656_),
    .Y(_15135_));
 sky130_fd_sc_hd__nand3_4 _37496_ (.A(_15107_),
    .B(_15134_),
    .C(_15135_),
    .Y(_15136_));
 sky130_fd_sc_hd__nand3_2 _37497_ (.A(_15129_),
    .B(_15133_),
    .C(_13663_),
    .Y(_15137_));
 sky130_fd_sc_hd__o2bb2ai_1 _37498_ (.A1_N(_15133_),
    .A2_N(_15129_),
    .B1(_13653_),
    .B2(_13651_),
    .Y(_15138_));
 sky130_fd_sc_hd__o211ai_4 _37499_ (.A1(_15106_),
    .A2(_14832_),
    .B1(_15137_),
    .C1(_15138_),
    .Y(_15139_));
 sky130_fd_sc_hd__o21ai_2 _37500_ (.A1(_13656_),
    .A2(_14863_),
    .B1(_14871_),
    .Y(_15140_));
 sky130_fd_sc_hd__a21oi_4 _37501_ (.A1(_15136_),
    .A2(_15139_),
    .B1(_15140_),
    .Y(_15141_));
 sky130_fd_sc_hd__nor2_1 _37502_ (.A(_14283_),
    .B(_14863_),
    .Y(_15142_));
 sky130_fd_sc_hd__o211a_4 _37503_ (.A1(_14864_),
    .A2(_15142_),
    .B1(_15139_),
    .C1(_15136_),
    .X(_15143_));
 sky130_fd_sc_hd__o2bb2ai_4 _37504_ (.A1_N(_15096_),
    .A2_N(_15105_),
    .B1(_15141_),
    .B2(_15143_),
    .Y(_15144_));
 sky130_fd_sc_hd__nor2_8 _37505_ (.A(_15141_),
    .B(_15143_),
    .Y(_15145_));
 sky130_fd_sc_hd__nand3_4 _37506_ (.A(_15105_),
    .B(_15096_),
    .C(_15145_),
    .Y(_15146_));
 sky130_fd_sc_hd__nand2_4 _37507_ (.A(_14894_),
    .B(_14835_),
    .Y(_15147_));
 sky130_fd_sc_hd__a21oi_4 _37508_ (.A1(_15144_),
    .A2(_15146_),
    .B1(_15147_),
    .Y(_15148_));
 sky130_fd_sc_hd__nand2_1 _37509_ (.A(_14831_),
    .B(_14834_),
    .Y(_15149_));
 sky130_fd_sc_hd__a21o_1 _37510_ (.A1(_14873_),
    .A2(_14878_),
    .B1(_14879_),
    .X(_15150_));
 sky130_fd_sc_hd__nand3_2 _37511_ (.A(_14873_),
    .B(_14878_),
    .C(_14879_),
    .Y(_15151_));
 sky130_fd_sc_hd__nand2_1 _37512_ (.A(_15150_),
    .B(_15151_),
    .Y(_15152_));
 sky130_fd_sc_hd__a21oi_1 _37513_ (.A1(_14836_),
    .A2(_15149_),
    .B1(_15152_),
    .Y(_15153_));
 sky130_fd_sc_hd__o211a_2 _37514_ (.A1(_14893_),
    .A2(_15153_),
    .B1(_15146_),
    .C1(_15144_),
    .X(_15154_));
 sky130_fd_sc_hd__nand2_2 _37515_ (.A(_15151_),
    .B(_14878_),
    .Y(_15155_));
 sky130_fd_sc_hd__nor2_4 _37516_ (.A(_14592_),
    .B(_15155_),
    .Y(_15156_));
 sky130_vsdinv _37517_ (.A(_15155_),
    .Y(_15157_));
 sky130_fd_sc_hd__nor2_8 _37518_ (.A(net411),
    .B(_15157_),
    .Y(_15158_));
 sky130_fd_sc_hd__nor2_4 _37519_ (.A(_15156_),
    .B(_15158_),
    .Y(_15159_));
 sky130_fd_sc_hd__o21ai_4 _37520_ (.A1(_15148_),
    .A2(_15154_),
    .B1(_15159_),
    .Y(_15160_));
 sky130_fd_sc_hd__o21a_2 _37521_ (.A1(_14899_),
    .A2(_14892_),
    .B1(_14898_),
    .X(_15161_));
 sky130_fd_sc_hd__a21o_1 _37522_ (.A1(_15144_),
    .A2(_15146_),
    .B1(_15147_),
    .X(_15162_));
 sky130_fd_sc_hd__nand3_4 _37523_ (.A(_15147_),
    .B(_15144_),
    .C(_15146_),
    .Y(_15163_));
 sky130_fd_sc_hd__nand2_1 _37524_ (.A(_15157_),
    .B(_14595_),
    .Y(_15164_));
 sky130_fd_sc_hd__or2b_4 _37525_ (.A(_15158_),
    .B_N(_15164_),
    .X(_15165_));
 sky130_fd_sc_hd__nand3_4 _37526_ (.A(_15162_),
    .B(_15163_),
    .C(_15165_),
    .Y(_15166_));
 sky130_fd_sc_hd__nand3_4 _37527_ (.A(_15160_),
    .B(_15161_),
    .C(_15166_),
    .Y(_15167_));
 sky130_fd_sc_hd__o22ai_4 _37528_ (.A1(_15158_),
    .A2(_15156_),
    .B1(_15148_),
    .B2(_15154_),
    .Y(_15168_));
 sky130_fd_sc_hd__o21ai_2 _37529_ (.A1(_14899_),
    .A2(_14892_),
    .B1(_14898_),
    .Y(_15169_));
 sky130_fd_sc_hd__nand3_4 _37530_ (.A(_15162_),
    .B(_15163_),
    .C(_15159_),
    .Y(_15170_));
 sky130_fd_sc_hd__nand3_4 _37531_ (.A(_15168_),
    .B(_15169_),
    .C(_15170_),
    .Y(_15171_));
 sky130_fd_sc_hd__a21oi_2 _37532_ (.A1(_15167_),
    .A2(_15171_),
    .B1(_14902_),
    .Y(_15172_));
 sky130_fd_sc_hd__and3_1 _37533_ (.A(_15167_),
    .B(_15171_),
    .C(_14902_),
    .X(_15173_));
 sky130_vsdinv _37534_ (.A(_14908_),
    .Y(_15174_));
 sky130_fd_sc_hd__nand2_1 _37535_ (.A(_14905_),
    .B(_14907_),
    .Y(_15175_));
 sky130_fd_sc_hd__a21boi_4 _37536_ (.A1(_15175_),
    .A2(_14631_),
    .B1_N(_14597_),
    .Y(_15176_));
 sky130_fd_sc_hd__nor2_2 _37537_ (.A(_15174_),
    .B(_15176_),
    .Y(_15177_));
 sky130_fd_sc_hd__o21ai_4 _37538_ (.A1(_15172_),
    .A2(_15173_),
    .B1(_15177_),
    .Y(_15178_));
 sky130_fd_sc_hd__nand3_2 _37539_ (.A(_15167_),
    .B(_15171_),
    .C(_14902_),
    .Y(_15179_));
 sky130_fd_sc_hd__nand2_1 _37540_ (.A(_15167_),
    .B(_15171_),
    .Y(_15180_));
 sky130_vsdinv _37541_ (.A(_14902_),
    .Y(_15181_));
 sky130_fd_sc_hd__nand2_1 _37542_ (.A(_15180_),
    .B(_15181_),
    .Y(_15182_));
 sky130_fd_sc_hd__o211ai_4 _37543_ (.A1(_15174_),
    .A2(_15176_),
    .B1(_15179_),
    .C1(_15182_),
    .Y(_15183_));
 sky130_fd_sc_hd__nand2_2 _37544_ (.A(_15178_),
    .B(_15183_),
    .Y(_15184_));
 sky130_fd_sc_hd__o2111a_1 _37545_ (.A1(_14910_),
    .A2(_14914_),
    .B1(_14626_),
    .C1(_14620_),
    .D1(_14915_),
    .X(_15185_));
 sky130_fd_sc_hd__o2111ai_4 _37546_ (.A1(_14910_),
    .A2(_14914_),
    .B1(_14626_),
    .C1(_14620_),
    .D1(_14915_),
    .Y(_15186_));
 sky130_fd_sc_hd__a21oi_1 _37547_ (.A1(_14911_),
    .A2(_14909_),
    .B1(_14913_),
    .Y(_15187_));
 sky130_fd_sc_hd__o22ai_1 _37548_ (.A1(_14910_),
    .A2(_14914_),
    .B1(_14626_),
    .B2(_15187_),
    .Y(_15188_));
 sky130_fd_sc_hd__o21bai_1 _37549_ (.A1(_15186_),
    .A2(_14629_),
    .B1_N(_15188_),
    .Y(_15189_));
 sky130_fd_sc_hd__a31o_4 _37550_ (.A1(_14034_),
    .A2(_14340_),
    .A3(_15185_),
    .B1(_15189_),
    .X(_15190_));
 sky130_fd_sc_hd__xnor2_4 _37551_ (.A(_15184_),
    .B(_15190_),
    .Y(_02663_));
 sky130_fd_sc_hd__and3_2 _37552_ (.A(_15168_),
    .B(_15169_),
    .C(_15170_),
    .X(_15191_));
 sky130_fd_sc_hd__a21oi_2 _37553_ (.A1(_15167_),
    .A2(_14902_),
    .B1(_15191_),
    .Y(_15192_));
 sky130_fd_sc_hd__a21bo_2 _37554_ (.A1(_15136_),
    .A2(_15140_),
    .B1_N(_15139_),
    .X(_15193_));
 sky130_fd_sc_hd__nor2_4 _37555_ (.A(_14305_),
    .B(_15193_),
    .Y(_15194_));
 sky130_fd_sc_hd__and2_1 _37556_ (.A(_15193_),
    .B(_13718_),
    .X(_15195_));
 sky130_fd_sc_hd__buf_2 _37557_ (.A(_15195_),
    .X(_15196_));
 sky130_fd_sc_hd__nor2_4 _37558_ (.A(_15194_),
    .B(_15196_),
    .Y(_15197_));
 sky130_fd_sc_hd__o21a_1 _37559_ (.A1(_14996_),
    .A2(_14985_),
    .B1(_15000_),
    .X(_15198_));
 sky130_fd_sc_hd__a21o_1 _37560_ (.A1(_14980_),
    .A2(_14982_),
    .B1(_14977_),
    .X(_15199_));
 sky130_fd_sc_hd__nand2_1 _37561_ (.A(_11079_),
    .B(_07330_),
    .Y(_15200_));
 sky130_fd_sc_hd__nand3b_4 _37562_ (.A_N(_15200_),
    .B(_12781_),
    .C(net440),
    .Y(_15201_));
 sky130_fd_sc_hd__o21ai_2 _37563_ (.A1(_06284_),
    .A2(_13099_),
    .B1(_15200_),
    .Y(_15202_));
 sky130_fd_sc_hd__nand2_2 _37564_ (.A(_10828_),
    .B(_07323_),
    .Y(_15203_));
 sky130_vsdinv _37565_ (.A(_15203_),
    .Y(_15204_));
 sky130_fd_sc_hd__a21o_1 _37566_ (.A1(_15201_),
    .A2(_15202_),
    .B1(_15204_),
    .X(_15205_));
 sky130_fd_sc_hd__nand3_2 _37567_ (.A(_15201_),
    .B(_15202_),
    .C(_15204_),
    .Y(_15206_));
 sky130_fd_sc_hd__nand3_4 _37568_ (.A(_15199_),
    .B(_15205_),
    .C(_15206_),
    .Y(_15207_));
 sky130_fd_sc_hd__a21oi_2 _37569_ (.A1(_15201_),
    .A2(_15202_),
    .B1(_15204_),
    .Y(_15208_));
 sky130_fd_sc_hd__o21a_1 _37570_ (.A1(_19892_),
    .A2(_13745_),
    .B1(_15200_),
    .X(_15209_));
 sky130_fd_sc_hd__a41o_1 _37571_ (.A1(_07275_),
    .A2(_12781_),
    .A3(_12779_),
    .A4(_11848_),
    .B1(_15203_),
    .X(_15210_));
 sky130_fd_sc_hd__nor2_2 _37572_ (.A(_15209_),
    .B(_15210_),
    .Y(_15211_));
 sky130_fd_sc_hd__a21oi_2 _37573_ (.A1(_14980_),
    .A2(_14982_),
    .B1(_14977_),
    .Y(_15212_));
 sky130_fd_sc_hd__o21ai_4 _37574_ (.A1(_15208_),
    .A2(_15211_),
    .B1(_15212_),
    .Y(_15213_));
 sky130_fd_sc_hd__nand2_4 _37575_ (.A(_11348_),
    .B(_06803_),
    .Y(_15214_));
 sky130_fd_sc_hd__nand2_4 _37576_ (.A(_10046_),
    .B(_06783_),
    .Y(_15215_));
 sky130_fd_sc_hd__nor2_4 _37577_ (.A(_15214_),
    .B(_15215_),
    .Y(_15216_));
 sky130_fd_sc_hd__and2_1 _37578_ (.A(_15214_),
    .B(_15215_),
    .X(_15217_));
 sky130_fd_sc_hd__nand2_1 _37579_ (.A(_19592_),
    .B(_10733_),
    .Y(_15218_));
 sky130_vsdinv _37580_ (.A(_15218_),
    .Y(_15219_));
 sky130_fd_sc_hd__o21ai_2 _37581_ (.A1(_15216_),
    .A2(_15217_),
    .B1(_15219_),
    .Y(_15220_));
 sky130_vsdinv _37582_ (.A(_15220_),
    .Y(_15221_));
 sky130_fd_sc_hd__nor2_1 _37583_ (.A(_15216_),
    .B(_15217_),
    .Y(_15222_));
 sky130_fd_sc_hd__nand2_2 _37584_ (.A(_15222_),
    .B(_15218_),
    .Y(_15223_));
 sky130_vsdinv _37585_ (.A(_15223_),
    .Y(_15224_));
 sky130_fd_sc_hd__o2bb2ai_1 _37586_ (.A1_N(_15207_),
    .A2_N(_15213_),
    .B1(_15221_),
    .B2(_15224_),
    .Y(_15225_));
 sky130_fd_sc_hd__nand2_4 _37587_ (.A(_15223_),
    .B(_15220_),
    .Y(_15226_));
 sky130_fd_sc_hd__nand3b_2 _37588_ (.A_N(_15226_),
    .B(_15213_),
    .C(_15207_),
    .Y(_15227_));
 sky130_fd_sc_hd__nand3_4 _37589_ (.A(_15198_),
    .B(_15225_),
    .C(_15227_),
    .Y(_15228_));
 sky130_fd_sc_hd__a21o_1 _37590_ (.A1(_15213_),
    .A2(_15207_),
    .B1(_15226_),
    .X(_15229_));
 sky130_fd_sc_hd__o21ai_2 _37591_ (.A1(_14996_),
    .A2(_14985_),
    .B1(_15000_),
    .Y(_15230_));
 sky130_fd_sc_hd__nand3_2 _37592_ (.A(_15213_),
    .B(_15207_),
    .C(_15226_),
    .Y(_15231_));
 sky130_fd_sc_hd__nand3_4 _37593_ (.A(_15229_),
    .B(_15230_),
    .C(_15231_),
    .Y(_15232_));
 sky130_fd_sc_hd__nand2_2 _37594_ (.A(_15228_),
    .B(_15232_),
    .Y(_15233_));
 sky130_fd_sc_hd__nor2_4 _37595_ (.A(_14989_),
    .B(_14992_),
    .Y(_15234_));
 sky130_fd_sc_hd__nor2_4 _37596_ (.A(_14993_),
    .B(_15234_),
    .Y(_15235_));
 sky130_fd_sc_hd__nand2_1 _37597_ (.A(_09485_),
    .B(_19871_),
    .Y(_15236_));
 sky130_fd_sc_hd__nand2_2 _37598_ (.A(_19600_),
    .B(_07705_),
    .Y(_15237_));
 sky130_fd_sc_hd__nor2_2 _37599_ (.A(_15236_),
    .B(_15237_),
    .Y(_15238_));
 sky130_fd_sc_hd__and2_1 _37600_ (.A(_15236_),
    .B(_15237_),
    .X(_15239_));
 sky130_fd_sc_hd__nor2_2 _37601_ (.A(_08579_),
    .B(_12916_),
    .Y(_15240_));
 sky130_fd_sc_hd__o21bai_4 _37602_ (.A1(_15238_),
    .A2(_15239_),
    .B1_N(_15240_),
    .Y(_15241_));
 sky130_vsdinv _37603_ (.A(_15238_),
    .Y(_15242_));
 sky130_fd_sc_hd__nand2_1 _37604_ (.A(_15236_),
    .B(_15237_),
    .Y(_15243_));
 sky130_fd_sc_hd__nand3_4 _37605_ (.A(_15242_),
    .B(_15240_),
    .C(_15243_),
    .Y(_15244_));
 sky130_fd_sc_hd__nand3_4 _37606_ (.A(_15235_),
    .B(_15241_),
    .C(_15244_),
    .Y(_15245_));
 sky130_fd_sc_hd__and2_2 _37607_ (.A(_15012_),
    .B(_15009_),
    .X(_15246_));
 sky130_fd_sc_hd__a21oi_4 _37608_ (.A1(_15244_),
    .A2(_15241_),
    .B1(_15235_),
    .Y(_15247_));
 sky130_fd_sc_hd__nor2_2 _37609_ (.A(_15246_),
    .B(_15247_),
    .Y(_15248_));
 sky130_fd_sc_hd__o2bb2ai_2 _37610_ (.A1_N(_15241_),
    .A2_N(_15244_),
    .B1(_14993_),
    .B2(_15234_),
    .Y(_15249_));
 sky130_fd_sc_hd__a21boi_4 _37611_ (.A1(_15249_),
    .A2(_15245_),
    .B1_N(_15246_),
    .Y(_15250_));
 sky130_fd_sc_hd__a21oi_4 _37612_ (.A1(_15245_),
    .A2(_15248_),
    .B1(_15250_),
    .Y(_15251_));
 sky130_fd_sc_hd__nand2_4 _37613_ (.A(_15233_),
    .B(_15251_),
    .Y(_15252_));
 sky130_fd_sc_hd__a21oi_4 _37614_ (.A1(_15003_),
    .A2(_15005_),
    .B1(_15004_),
    .Y(_15253_));
 sky130_fd_sc_hd__a21oi_4 _37615_ (.A1(_15006_),
    .A2(_15031_),
    .B1(_15253_),
    .Y(_15254_));
 sky130_fd_sc_hd__a21o_1 _37616_ (.A1(_15245_),
    .A2(_15248_),
    .B1(_15250_),
    .X(_15255_));
 sky130_fd_sc_hd__nand3_4 _37617_ (.A(_15255_),
    .B(_15228_),
    .C(_15232_),
    .Y(_15256_));
 sky130_fd_sc_hd__nand3_4 _37618_ (.A(_15252_),
    .B(_15254_),
    .C(_15256_),
    .Y(_15257_));
 sky130_fd_sc_hd__a31oi_4 _37619_ (.A1(_15004_),
    .A2(_15005_),
    .A3(_15003_),
    .B1(_15039_),
    .Y(_15258_));
 sky130_fd_sc_hd__nand3_2 _37620_ (.A(_15251_),
    .B(_15228_),
    .C(_15232_),
    .Y(_15259_));
 sky130_fd_sc_hd__nand2_1 _37621_ (.A(_15233_),
    .B(_15255_),
    .Y(_15260_));
 sky130_fd_sc_hd__o211ai_4 _37622_ (.A1(_15253_),
    .A2(_15258_),
    .B1(_15259_),
    .C1(_15260_),
    .Y(_15261_));
 sky130_fd_sc_hd__a22oi_4 _37623_ (.A1(_11847_),
    .A2(_09823_),
    .B1(_11849_),
    .B2(_11909_),
    .Y(_15262_));
 sky130_fd_sc_hd__and4_2 _37624_ (.A(_07934_),
    .B(_07758_),
    .C(_19848_),
    .D(_09075_),
    .X(_15263_));
 sky130_fd_sc_hd__a211o_1 _37625_ (.A1(_13408_),
    .A2(_13248_),
    .B1(_15262_),
    .C1(_15263_),
    .X(_15264_));
 sky130_fd_sc_hd__nor2_1 _37626_ (.A(net471),
    .B(_13900_),
    .Y(_15265_));
 sky130_fd_sc_hd__o21ai_2 _37627_ (.A1(_15262_),
    .A2(_15263_),
    .B1(_15265_),
    .Y(_15266_));
 sky130_fd_sc_hd__nand2_4 _37628_ (.A(_15264_),
    .B(_15266_),
    .Y(_15267_));
 sky130_fd_sc_hd__nand2_2 _37629_ (.A(_08153_),
    .B(_10458_),
    .Y(_15268_));
 sky130_fd_sc_hd__nand2_2 _37630_ (.A(_08155_),
    .B(_10453_),
    .Y(_15269_));
 sky130_fd_sc_hd__nor2_4 _37631_ (.A(_15268_),
    .B(_15269_),
    .Y(_15270_));
 sky130_fd_sc_hd__and2_1 _37632_ (.A(_15268_),
    .B(_15269_),
    .X(_15271_));
 sky130_fd_sc_hd__nand2_2 _37633_ (.A(_19617_),
    .B(_11232_),
    .Y(_15272_));
 sky130_fd_sc_hd__o21ai_2 _37634_ (.A1(_15270_),
    .A2(_15271_),
    .B1(_15272_),
    .Y(_15273_));
 sky130_fd_sc_hd__or2_1 _37635_ (.A(_15268_),
    .B(_15269_),
    .X(_15274_));
 sky130_fd_sc_hd__nand2_2 _37636_ (.A(_15268_),
    .B(_15269_),
    .Y(_15275_));
 sky130_vsdinv _37637_ (.A(_15272_),
    .Y(_15276_));
 sky130_fd_sc_hd__nand3_2 _37638_ (.A(_15274_),
    .B(_15275_),
    .C(_15276_),
    .Y(_15277_));
 sky130_fd_sc_hd__a21o_1 _37639_ (.A1(_15050_),
    .A2(_15049_),
    .B1(_15045_),
    .X(_15278_));
 sky130_fd_sc_hd__nand3_4 _37640_ (.A(_15273_),
    .B(_15277_),
    .C(_15278_),
    .Y(_15279_));
 sky130_fd_sc_hd__o21ai_2 _37641_ (.A1(_15270_),
    .A2(_15271_),
    .B1(_15276_),
    .Y(_15280_));
 sky130_fd_sc_hd__nand3_2 _37642_ (.A(_15274_),
    .B(_15275_),
    .C(_15272_),
    .Y(_15281_));
 sky130_fd_sc_hd__a21oi_2 _37643_ (.A1(_15050_),
    .A2(_15049_),
    .B1(_15045_),
    .Y(_15282_));
 sky130_fd_sc_hd__nand3_4 _37644_ (.A(_15280_),
    .B(_15281_),
    .C(_15282_),
    .Y(_15283_));
 sky130_fd_sc_hd__nand3_4 _37645_ (.A(_15267_),
    .B(_15279_),
    .C(_15283_),
    .Y(_15284_));
 sky130_fd_sc_hd__a21o_2 _37646_ (.A1(_15279_),
    .A2(_15283_),
    .B1(_15267_),
    .X(_15285_));
 sky130_fd_sc_hd__nor2_2 _37647_ (.A(_15021_),
    .B(_15024_),
    .Y(_15286_));
 sky130_fd_sc_hd__o2bb2ai_4 _37648_ (.A1_N(_15284_),
    .A2_N(_15285_),
    .B1(_15036_),
    .B2(_15286_),
    .Y(_15287_));
 sky130_fd_sc_hd__o21ai_2 _37649_ (.A1(_15036_),
    .A2(_15037_),
    .B1(_15020_),
    .Y(_15288_));
 sky130_fd_sc_hd__nand3_4 _37650_ (.A(_15288_),
    .B(_15285_),
    .C(_15284_),
    .Y(_15289_));
 sky130_fd_sc_hd__nand2_2 _37651_ (.A(_15069_),
    .B(_15057_),
    .Y(_15290_));
 sky130_fd_sc_hd__nand2_4 _37652_ (.A(_15290_),
    .B(_15053_),
    .Y(_15291_));
 sky130_fd_sc_hd__a21oi_4 _37653_ (.A1(_15287_),
    .A2(_15289_),
    .B1(_15291_),
    .Y(_15292_));
 sky130_fd_sc_hd__and3_1 _37654_ (.A(_15287_),
    .B(_15289_),
    .C(_15291_),
    .X(_15293_));
 sky130_fd_sc_hd__o2bb2ai_4 _37655_ (.A1_N(_15257_),
    .A2_N(_15261_),
    .B1(_15292_),
    .B2(_15293_),
    .Y(_15294_));
 sky130_fd_sc_hd__nor2_2 _37656_ (.A(_15292_),
    .B(_15293_),
    .Y(_15295_));
 sky130_fd_sc_hd__nand3_4 _37657_ (.A(_15295_),
    .B(_15261_),
    .C(_15257_),
    .Y(_15296_));
 sky130_fd_sc_hd__nand2_1 _37658_ (.A(_15082_),
    .B(_15042_),
    .Y(_15297_));
 sky130_fd_sc_hd__nand2_4 _37659_ (.A(_15297_),
    .B(_15033_),
    .Y(_15298_));
 sky130_fd_sc_hd__a21oi_4 _37660_ (.A1(_15294_),
    .A2(_15296_),
    .B1(_15298_),
    .Y(_15299_));
 sky130_vsdinv _37661_ (.A(_15033_),
    .Y(_15300_));
 sky130_vsdinv _37662_ (.A(_15053_),
    .Y(_15301_));
 sky130_fd_sc_hd__o211a_1 _37663_ (.A1(_15301_),
    .A2(_15290_),
    .B1(_15068_),
    .C1(_15071_),
    .X(_15302_));
 sky130_fd_sc_hd__o21ai_1 _37664_ (.A1(_15079_),
    .A2(_15302_),
    .B1(_15080_),
    .Y(_15303_));
 sky130_fd_sc_hd__nand2_1 _37665_ (.A(_15303_),
    .B(_15076_),
    .Y(_15304_));
 sky130_fd_sc_hd__a31oi_1 _37666_ (.A1(_15041_),
    .A2(_15040_),
    .A3(_15035_),
    .B1(_15304_),
    .Y(_15305_));
 sky130_fd_sc_hd__o211a_2 _37667_ (.A1(_15300_),
    .A2(_15305_),
    .B1(_15296_),
    .C1(_15294_),
    .X(_15306_));
 sky130_fd_sc_hd__nand2_1 _37668_ (.A(_11695_),
    .B(_10488_),
    .Y(_15307_));
 sky130_fd_sc_hd__nand2_1 _37669_ (.A(_08873_),
    .B(_09933_),
    .Y(_15308_));
 sky130_fd_sc_hd__or2_2 _37670_ (.A(_15307_),
    .B(_15308_),
    .X(_15309_));
 sky130_fd_sc_hd__nor2_2 _37671_ (.A(net441),
    .B(_10596_),
    .Y(_15310_));
 sky130_fd_sc_hd__nand2_1 _37672_ (.A(_15307_),
    .B(_15308_),
    .Y(_15311_));
 sky130_fd_sc_hd__nand3_4 _37673_ (.A(_15309_),
    .B(_15310_),
    .C(_15311_),
    .Y(_15312_));
 sky130_fd_sc_hd__a21o_1 _37674_ (.A1(_10991_),
    .A2(_12639_),
    .B1(_15307_),
    .X(_15313_));
 sky130_fd_sc_hd__a21o_1 _37675_ (.A1(_10990_),
    .A2(_11179_),
    .B1(_15308_),
    .X(_15314_));
 sky130_fd_sc_hd__nand3b_4 _37676_ (.A_N(_15310_),
    .B(_15313_),
    .C(_15314_),
    .Y(_15315_));
 sky130_fd_sc_hd__clkbuf_4 _37677_ (.A(_09359_),
    .X(_15316_));
 sky130_fd_sc_hd__a31o_2 _37678_ (.A1(_15062_),
    .A2(_13408_),
    .A3(_15316_),
    .B1(_15061_),
    .X(_15317_));
 sky130_fd_sc_hd__a21oi_2 _37679_ (.A1(_15312_),
    .A2(_15315_),
    .B1(_15317_),
    .Y(_15318_));
 sky130_fd_sc_hd__a21oi_1 _37680_ (.A1(_15059_),
    .A2(_15060_),
    .B1(_15064_),
    .Y(_15319_));
 sky130_fd_sc_hd__o211a_1 _37681_ (.A1(_15061_),
    .A2(_15319_),
    .B1(_15315_),
    .C1(_15312_),
    .X(_15320_));
 sky130_fd_sc_hd__nand2_2 _37682_ (.A(_14926_),
    .B(_14924_),
    .Y(_15321_));
 sky130_fd_sc_hd__o21bai_4 _37683_ (.A1(_15318_),
    .A2(_15320_),
    .B1_N(_15321_),
    .Y(_15322_));
 sky130_fd_sc_hd__a21o_1 _37684_ (.A1(_15312_),
    .A2(_15315_),
    .B1(_15317_),
    .X(_15323_));
 sky130_fd_sc_hd__nand3_4 _37685_ (.A(_15312_),
    .B(_15317_),
    .C(_15315_),
    .Y(_15324_));
 sky130_fd_sc_hd__nand3_4 _37686_ (.A(_15323_),
    .B(_15321_),
    .C(_15324_),
    .Y(_15325_));
 sky130_fd_sc_hd__o21ai_4 _37687_ (.A1(_14933_),
    .A2(_14929_),
    .B1(_14936_),
    .Y(_15326_));
 sky130_fd_sc_hd__a21oi_4 _37688_ (.A1(_15322_),
    .A2(_15325_),
    .B1(_15326_),
    .Y(_15327_));
 sky130_fd_sc_hd__nand2_2 _37689_ (.A(_15323_),
    .B(_15321_),
    .Y(_15328_));
 sky130_fd_sc_hd__o211a_1 _37690_ (.A1(_15320_),
    .A2(_15328_),
    .B1(_15322_),
    .C1(_15326_),
    .X(_15329_));
 sky130_fd_sc_hd__nand2_2 _37691_ (.A(_19644_),
    .B(_10613_),
    .Y(_15330_));
 sky130_fd_sc_hd__nand2_2 _37692_ (.A(_11593_),
    .B(_06416_),
    .Y(_15331_));
 sky130_fd_sc_hd__o21ai_1 _37693_ (.A1(_15330_),
    .A2(_15331_),
    .B1(_14946_),
    .Y(_15332_));
 sky130_fd_sc_hd__a21o_1 _37694_ (.A1(_15330_),
    .A2(_15331_),
    .B1(_15332_),
    .X(_15333_));
 sky130_fd_sc_hd__nor2_1 _37695_ (.A(_15330_),
    .B(_15331_),
    .Y(_15334_));
 sky130_fd_sc_hd__and2_1 _37696_ (.A(_15330_),
    .B(_15331_),
    .X(_15335_));
 sky130_fd_sc_hd__o21ai_2 _37697_ (.A1(_15334_),
    .A2(_15335_),
    .B1(_14947_),
    .Y(_15336_));
 sky130_fd_sc_hd__a21oi_4 _37698_ (.A1(_14947_),
    .A2(_14948_),
    .B1(_14945_),
    .Y(_15337_));
 sky130_fd_sc_hd__nand3_4 _37699_ (.A(_15333_),
    .B(_15336_),
    .C(_15337_),
    .Y(_15338_));
 sky130_fd_sc_hd__a21o_2 _37700_ (.A1(_15333_),
    .A2(_15336_),
    .B1(_15337_),
    .X(_15339_));
 sky130_fd_sc_hd__o2bb2ai_2 _37701_ (.A1_N(_15338_),
    .A2_N(_15339_),
    .B1(_14807_),
    .B2(_14803_),
    .Y(_15340_));
 sky130_fd_sc_hd__nand3_4 _37702_ (.A(_15339_),
    .B(_14809_),
    .C(_15338_),
    .Y(_15341_));
 sky130_fd_sc_hd__nand2_2 _37703_ (.A(_15340_),
    .B(_15341_),
    .Y(_15342_));
 sky130_fd_sc_hd__o21ai_2 _37704_ (.A1(_15327_),
    .A2(_15329_),
    .B1(_15342_),
    .Y(_15343_));
 sky130_fd_sc_hd__nor2_2 _37705_ (.A(_14937_),
    .B(_14932_),
    .Y(_15344_));
 sky130_fd_sc_hd__o2bb2ai_4 _37706_ (.A1_N(_15322_),
    .A2_N(_15325_),
    .B1(_14929_),
    .B2(_15344_),
    .Y(_15345_));
 sky130_fd_sc_hd__nand3_4 _37707_ (.A(_15326_),
    .B(_15322_),
    .C(_15325_),
    .Y(_15346_));
 sky130_fd_sc_hd__nand3b_4 _37708_ (.A_N(_15342_),
    .B(_15345_),
    .C(_15346_),
    .Y(_15347_));
 sky130_fd_sc_hd__o21ai_4 _37709_ (.A1(_15079_),
    .A2(_15080_),
    .B1(_15073_),
    .Y(_15348_));
 sky130_fd_sc_hd__a21oi_1 _37710_ (.A1(_15343_),
    .A2(_15347_),
    .B1(_15348_),
    .Y(_15349_));
 sky130_fd_sc_hd__o211a_1 _37711_ (.A1(_15302_),
    .A2(_15081_),
    .B1(_15347_),
    .C1(_15343_),
    .X(_15350_));
 sky130_fd_sc_hd__o21ai_4 _37712_ (.A1(_14940_),
    .A2(_14965_),
    .B1(_14964_),
    .Y(_15351_));
 sky130_vsdinv _37713_ (.A(_15351_),
    .Y(_15352_));
 sky130_fd_sc_hd__o21ai_1 _37714_ (.A1(_15349_),
    .A2(_15350_),
    .B1(_15352_),
    .Y(_15353_));
 sky130_fd_sc_hd__a22oi_4 _37715_ (.A1(_15340_),
    .A2(_15341_),
    .B1(_15345_),
    .B2(_15346_),
    .Y(_15354_));
 sky130_fd_sc_hd__nor3_4 _37716_ (.A(_15342_),
    .B(_15327_),
    .C(_15329_),
    .Y(_15355_));
 sky130_fd_sc_hd__o21bai_4 _37717_ (.A1(_15354_),
    .A2(_15355_),
    .B1_N(_15348_),
    .Y(_15356_));
 sky130_fd_sc_hd__nand3_4 _37718_ (.A(_15343_),
    .B(_15348_),
    .C(_15347_),
    .Y(_15357_));
 sky130_fd_sc_hd__nand3_1 _37719_ (.A(_15356_),
    .B(_15357_),
    .C(_15351_),
    .Y(_15358_));
 sky130_fd_sc_hd__nand2_2 _37720_ (.A(_15353_),
    .B(_15358_),
    .Y(_15359_));
 sky130_fd_sc_hd__o21bai_2 _37721_ (.A1(_15299_),
    .A2(_15306_),
    .B1_N(_15359_),
    .Y(_15360_));
 sky130_fd_sc_hd__nand2_1 _37722_ (.A(_15101_),
    .B(_15092_),
    .Y(_15361_));
 sky130_fd_sc_hd__nand2_1 _37723_ (.A(_15361_),
    .B(_15090_),
    .Y(_15362_));
 sky130_fd_sc_hd__a21o_1 _37724_ (.A1(_15294_),
    .A2(_15296_),
    .B1(_15298_),
    .X(_15363_));
 sky130_fd_sc_hd__nand3_4 _37725_ (.A(_15298_),
    .B(_15294_),
    .C(_15296_),
    .Y(_15364_));
 sky130_fd_sc_hd__nand3_2 _37726_ (.A(_15363_),
    .B(_15364_),
    .C(_15359_),
    .Y(_15365_));
 sky130_fd_sc_hd__nand3_4 _37727_ (.A(_15360_),
    .B(_15362_),
    .C(_15365_),
    .Y(_15366_));
 sky130_fd_sc_hd__a21oi_4 _37728_ (.A1(_15356_),
    .A2(_15357_),
    .B1(_15351_),
    .Y(_15367_));
 sky130_fd_sc_hd__nor2_1 _37729_ (.A(_14940_),
    .B(_14965_),
    .Y(_15368_));
 sky130_fd_sc_hd__o211a_1 _37730_ (.A1(_14942_),
    .A2(_15368_),
    .B1(_15357_),
    .C1(_15356_),
    .X(_15369_));
 sky130_fd_sc_hd__o22ai_4 _37731_ (.A1(_15367_),
    .A2(_15369_),
    .B1(_15299_),
    .B2(_15306_),
    .Y(_15370_));
 sky130_fd_sc_hd__nor2_2 _37732_ (.A(_15367_),
    .B(_15369_),
    .Y(_15371_));
 sky130_fd_sc_hd__nand3_4 _37733_ (.A(_15363_),
    .B(_15371_),
    .C(_15364_),
    .Y(_15372_));
 sky130_fd_sc_hd__o21ai_2 _37734_ (.A1(_15101_),
    .A2(_15086_),
    .B1(_15092_),
    .Y(_15373_));
 sky130_fd_sc_hd__nand3_4 _37735_ (.A(_15370_),
    .B(_15372_),
    .C(_15373_),
    .Y(_15374_));
 sky130_fd_sc_hd__nand2_1 _37736_ (.A(_15366_),
    .B(_15374_),
    .Y(_15375_));
 sky130_fd_sc_hd__nand3_4 _37737_ (.A(_15115_),
    .B(_14955_),
    .C(_14957_),
    .Y(_15376_));
 sky130_fd_sc_hd__a21oi_1 _37738_ (.A1(_14949_),
    .A2(_14952_),
    .B1(_14953_),
    .Y(_15377_));
 sky130_fd_sc_hd__o21ai_2 _37739_ (.A1(_14815_),
    .A2(_15377_),
    .B1(_14955_),
    .Y(_15378_));
 sky130_fd_sc_hd__nand3_4 _37740_ (.A(_15378_),
    .B(_15114_),
    .C(_15113_),
    .Y(_15379_));
 sky130_fd_sc_hd__nand2_2 _37741_ (.A(_15111_),
    .B(_14257_),
    .Y(_15380_));
 sky130_fd_sc_hd__nand2_4 _37742_ (.A(_15380_),
    .B(_15109_),
    .Y(_15381_));
 sky130_fd_sc_hd__a21oi_2 _37743_ (.A1(_15376_),
    .A2(_15379_),
    .B1(_15381_),
    .Y(_15382_));
 sky130_vsdinv _37744_ (.A(_15109_),
    .Y(_15383_));
 sky130_vsdinv _37745_ (.A(_15380_),
    .Y(_15384_));
 sky130_fd_sc_hd__o211a_1 _37746_ (.A1(_15383_),
    .A2(_15384_),
    .B1(_15379_),
    .C1(_15376_),
    .X(_15385_));
 sky130_fd_sc_hd__nor2_4 _37747_ (.A(_15116_),
    .B(_15115_),
    .Y(_15386_));
 sky130_fd_sc_hd__a2bb2oi_4 _37748_ (.A1_N(_15122_),
    .A2_N(_15123_),
    .B1(_15116_),
    .B2(_15115_),
    .Y(_15387_));
 sky130_fd_sc_hd__nor2_2 _37749_ (.A(_15386_),
    .B(_15387_),
    .Y(_15388_));
 sky130_fd_sc_hd__o21ai_4 _37750_ (.A1(_15382_),
    .A2(_15385_),
    .B1(_15388_),
    .Y(_15389_));
 sky130_fd_sc_hd__nand3_4 _37751_ (.A(_15376_),
    .B(_15379_),
    .C(_15381_),
    .Y(_15390_));
 sky130_fd_sc_hd__nand2_1 _37752_ (.A(_15376_),
    .B(_15379_),
    .Y(_15391_));
 sky130_vsdinv _37753_ (.A(_15381_),
    .Y(_15392_));
 sky130_fd_sc_hd__nand2_1 _37754_ (.A(_15391_),
    .B(_15392_),
    .Y(_15393_));
 sky130_fd_sc_hd__o211ai_4 _37755_ (.A1(_15386_),
    .A2(_15387_),
    .B1(_15390_),
    .C1(_15393_),
    .Y(_15394_));
 sky130_fd_sc_hd__a22oi_4 _37756_ (.A1(_13717_),
    .A2(_13939_),
    .B1(_15389_),
    .B2(_15394_),
    .Y(_15395_));
 sky130_fd_sc_hd__o2bb2ai_1 _37757_ (.A1_N(_15391_),
    .A2_N(_15392_),
    .B1(_15386_),
    .B2(_15387_),
    .Y(_15396_));
 sky130_fd_sc_hd__o211a_1 _37758_ (.A1(_15385_),
    .A2(_15396_),
    .B1(_13978_),
    .C1(_15389_),
    .X(_15397_));
 sky130_fd_sc_hd__a31oi_4 _37759_ (.A1(_14960_),
    .A2(_14962_),
    .A3(_14966_),
    .B1(_14972_),
    .Y(_15398_));
 sky130_fd_sc_hd__nor2_2 _37760_ (.A(_15097_),
    .B(_15398_),
    .Y(_15399_));
 sky130_fd_sc_hd__o21ai_4 _37761_ (.A1(_15395_),
    .A2(_15397_),
    .B1(_15399_),
    .Y(_15400_));
 sky130_fd_sc_hd__nand3_2 _37762_ (.A(_15389_),
    .B(_13988_),
    .C(_15394_),
    .Y(_15401_));
 sky130_fd_sc_hd__a21o_1 _37763_ (.A1(_15389_),
    .A2(_15394_),
    .B1(_13663_),
    .X(_15402_));
 sky130_fd_sc_hd__o211ai_4 _37764_ (.A1(_15097_),
    .A2(_15398_),
    .B1(_15401_),
    .C1(_15402_),
    .Y(_15403_));
 sky130_vsdinv _37765_ (.A(_15133_),
    .Y(_15404_));
 sky130_fd_sc_hd__a21o_1 _37766_ (.A1(_13989_),
    .A2(_15129_),
    .B1(_15404_),
    .X(_15405_));
 sky130_fd_sc_hd__a21oi_4 _37767_ (.A1(_15400_),
    .A2(_15403_),
    .B1(_15405_),
    .Y(_15406_));
 sky130_fd_sc_hd__and2_1 _37768_ (.A(_15129_),
    .B(_13988_),
    .X(_15407_));
 sky130_fd_sc_hd__o211a_4 _37769_ (.A1(_15404_),
    .A2(_15407_),
    .B1(_15403_),
    .C1(_15400_),
    .X(_15408_));
 sky130_fd_sc_hd__nor2_8 _37770_ (.A(_15406_),
    .B(_15408_),
    .Y(_15409_));
 sky130_fd_sc_hd__nand2_1 _37771_ (.A(_15375_),
    .B(_15409_),
    .Y(_15410_));
 sky130_fd_sc_hd__a21boi_4 _37772_ (.A1(_15105_),
    .A2(_15145_),
    .B1_N(_15096_),
    .Y(_15411_));
 sky130_fd_sc_hd__o211ai_4 _37773_ (.A1(_15406_),
    .A2(_15408_),
    .B1(_15374_),
    .C1(_15366_),
    .Y(_15412_));
 sky130_fd_sc_hd__nand3_4 _37774_ (.A(_15410_),
    .B(_15411_),
    .C(_15412_),
    .Y(_15413_));
 sky130_fd_sc_hd__o2bb2ai_1 _37775_ (.A1_N(_15366_),
    .A2_N(_15374_),
    .B1(_15406_),
    .B2(_15408_),
    .Y(_15414_));
 sky130_vsdinv _37776_ (.A(_15093_),
    .Y(_15415_));
 sky130_fd_sc_hd__nand2_1 _37777_ (.A(_15089_),
    .B(_15095_),
    .Y(_15416_));
 sky130_fd_sc_hd__o2bb2ai_2 _37778_ (.A1_N(_15145_),
    .A2_N(_15105_),
    .B1(_15415_),
    .B2(_15416_),
    .Y(_15417_));
 sky130_fd_sc_hd__nand3_2 _37779_ (.A(_15409_),
    .B(_15366_),
    .C(_15374_),
    .Y(_15418_));
 sky130_fd_sc_hd__nand3_4 _37780_ (.A(_15414_),
    .B(_15417_),
    .C(_15418_),
    .Y(_15419_));
 sky130_fd_sc_hd__nand3b_2 _37781_ (.A_N(_15197_),
    .B(_15413_),
    .C(_15419_),
    .Y(_15420_));
 sky130_fd_sc_hd__and2_1 _37782_ (.A(_15193_),
    .B(_14595_),
    .X(_15421_));
 sky130_fd_sc_hd__nor2_1 _37783_ (.A(_14329_),
    .B(_15193_),
    .Y(_15422_));
 sky130_fd_sc_hd__o2bb2ai_1 _37784_ (.A1_N(_15419_),
    .A2_N(_15413_),
    .B1(_15421_),
    .B2(_15422_),
    .Y(_15423_));
 sky130_fd_sc_hd__o2111ai_4 _37785_ (.A1(_15148_),
    .A2(_15165_),
    .B1(_15163_),
    .C1(_15420_),
    .D1(_15423_),
    .Y(_15424_));
 sky130_fd_sc_hd__o21ai_2 _37786_ (.A1(_15165_),
    .A2(_15148_),
    .B1(_15163_),
    .Y(_15425_));
 sky130_fd_sc_hd__o2bb2ai_2 _37787_ (.A1_N(_15419_),
    .A2_N(_15413_),
    .B1(_15196_),
    .B2(_15194_),
    .Y(_15426_));
 sky130_fd_sc_hd__nand3_4 _37788_ (.A(_15413_),
    .B(_15419_),
    .C(_15197_),
    .Y(_15427_));
 sky130_fd_sc_hd__nand3_4 _37789_ (.A(_15425_),
    .B(_15426_),
    .C(_15427_),
    .Y(_15428_));
 sky130_fd_sc_hd__nand2_1 _37790_ (.A(_15424_),
    .B(_15428_),
    .Y(_15429_));
 sky130_fd_sc_hd__nand2_1 _37791_ (.A(_15429_),
    .B(_15158_),
    .Y(_15430_));
 sky130_vsdinv _37792_ (.A(_15158_),
    .Y(_15431_));
 sky130_fd_sc_hd__nand3_2 _37793_ (.A(_15424_),
    .B(_15428_),
    .C(_15431_),
    .Y(_15432_));
 sky130_fd_sc_hd__nand3_4 _37794_ (.A(_15192_),
    .B(_15430_),
    .C(_15432_),
    .Y(_15433_));
 sky130_fd_sc_hd__a31oi_4 _37795_ (.A1(_15160_),
    .A2(_15161_),
    .A3(_15166_),
    .B1(_15181_),
    .Y(_15434_));
 sky130_fd_sc_hd__nand3_4 _37796_ (.A(_15424_),
    .B(_15428_),
    .C(_15158_),
    .Y(_15435_));
 sky130_fd_sc_hd__o2bb2ai_2 _37797_ (.A1_N(_15428_),
    .A2_N(_15424_),
    .B1(_14332_),
    .B2(_15157_),
    .Y(_15436_));
 sky130_fd_sc_hd__o211ai_4 _37798_ (.A1(_15191_),
    .A2(_15434_),
    .B1(_15435_),
    .C1(_15436_),
    .Y(_15437_));
 sky130_fd_sc_hd__nand2_2 _37799_ (.A(_15433_),
    .B(_15437_),
    .Y(_15438_));
 sky130_vsdinv _37800_ (.A(_15183_),
    .Y(_15439_));
 sky130_fd_sc_hd__a21oi_4 _37801_ (.A1(_15190_),
    .A2(_15178_),
    .B1(_15439_),
    .Y(_15440_));
 sky130_fd_sc_hd__xor2_4 _37802_ (.A(_15438_),
    .B(_15440_),
    .X(_02664_));
 sky130_fd_sc_hd__nand2_2 _37803_ (.A(_11695_),
    .B(_09933_),
    .Y(_15441_));
 sky130_fd_sc_hd__nand2_2 _37804_ (.A(_08623_),
    .B(_19829_),
    .Y(_15442_));
 sky130_fd_sc_hd__nor2_2 _37805_ (.A(_15441_),
    .B(_15442_),
    .Y(_15443_));
 sky130_fd_sc_hd__and2_1 _37806_ (.A(_15441_),
    .B(_15442_),
    .X(_15444_));
 sky130_fd_sc_hd__nor2_2 _37807_ (.A(net441),
    .B(_12618_),
    .Y(_15445_));
 sky130_fd_sc_hd__o21bai_4 _37808_ (.A1(_15443_),
    .A2(_15444_),
    .B1_N(_15445_),
    .Y(_15446_));
 sky130_fd_sc_hd__or2_2 _37809_ (.A(_15441_),
    .B(_15442_),
    .X(_15447_));
 sky130_fd_sc_hd__nand2_1 _37810_ (.A(_15441_),
    .B(_15442_),
    .Y(_15448_));
 sky130_fd_sc_hd__nand3_4 _37811_ (.A(_15447_),
    .B(_15445_),
    .C(_15448_),
    .Y(_15449_));
 sky130_fd_sc_hd__nand2_1 _37812_ (.A(_19628_),
    .B(_10493_),
    .Y(_15450_));
 sky130_fd_sc_hd__o21bai_4 _37813_ (.A1(_15450_),
    .A2(_15262_),
    .B1_N(_15263_),
    .Y(_15451_));
 sky130_fd_sc_hd__a21oi_4 _37814_ (.A1(_15446_),
    .A2(_15449_),
    .B1(_15451_),
    .Y(_15452_));
 sky130_fd_sc_hd__and3_2 _37815_ (.A(_15446_),
    .B(_15449_),
    .C(_15451_),
    .X(_15453_));
 sky130_fd_sc_hd__nand2_4 _37816_ (.A(_15312_),
    .B(_15309_),
    .Y(_15454_));
 sky130_vsdinv _37817_ (.A(_15454_),
    .Y(_15455_));
 sky130_fd_sc_hd__o21ai_4 _37818_ (.A1(_15452_),
    .A2(_15453_),
    .B1(_15455_),
    .Y(_15456_));
 sky130_fd_sc_hd__a21o_1 _37819_ (.A1(_15446_),
    .A2(_15449_),
    .B1(_15451_),
    .X(_15457_));
 sky130_fd_sc_hd__nand3_4 _37820_ (.A(_15446_),
    .B(_15449_),
    .C(_15451_),
    .Y(_15458_));
 sky130_fd_sc_hd__nand3_4 _37821_ (.A(_15457_),
    .B(_15454_),
    .C(_15458_),
    .Y(_15459_));
 sky130_fd_sc_hd__nand2_4 _37822_ (.A(_15328_),
    .B(_15324_),
    .Y(_15460_));
 sky130_fd_sc_hd__a21oi_4 _37823_ (.A1(_15456_),
    .A2(_15459_),
    .B1(_15460_),
    .Y(_15461_));
 sky130_fd_sc_hd__nand2_2 _37824_ (.A(_15457_),
    .B(_15454_),
    .Y(_15462_));
 sky130_fd_sc_hd__o211a_1 _37825_ (.A1(_15453_),
    .A2(_15462_),
    .B1(_15456_),
    .C1(_15460_),
    .X(_15463_));
 sky130_fd_sc_hd__o21ai_2 _37826_ (.A1(net445),
    .A2(_06423_),
    .B1(_11596_),
    .Y(_15464_));
 sky130_fd_sc_hd__and3_2 _37827_ (.A(_11184_),
    .B(_08219_),
    .C(_06168_),
    .X(_15465_));
 sky130_fd_sc_hd__nor2_1 _37828_ (.A(_15464_),
    .B(_15465_),
    .Y(_15466_));
 sky130_fd_sc_hd__o21ai_1 _37829_ (.A1(net473),
    .A2(_15335_),
    .B1(_15332_),
    .Y(_15467_));
 sky130_fd_sc_hd__or2_2 _37830_ (.A(_15466_),
    .B(_15467_),
    .X(_15468_));
 sky130_fd_sc_hd__nand2_2 _37831_ (.A(_15467_),
    .B(_15466_),
    .Y(_15469_));
 sky130_fd_sc_hd__nand2_2 _37832_ (.A(_15468_),
    .B(_15469_),
    .Y(_15470_));
 sky130_fd_sc_hd__nand2_2 _37833_ (.A(_15470_),
    .B(_14809_),
    .Y(_15471_));
 sky130_fd_sc_hd__nand3_4 _37834_ (.A(_15468_),
    .B(_14815_),
    .C(_15469_),
    .Y(_15472_));
 sky130_fd_sc_hd__nand2_2 _37835_ (.A(_15471_),
    .B(_15472_),
    .Y(_15473_));
 sky130_fd_sc_hd__o21ai_2 _37836_ (.A1(_15461_),
    .A2(_15463_),
    .B1(_15473_),
    .Y(_15474_));
 sky130_fd_sc_hd__nand3_2 _37837_ (.A(_15287_),
    .B(_15289_),
    .C(_15291_),
    .Y(_15475_));
 sky130_fd_sc_hd__nand2_2 _37838_ (.A(_15475_),
    .B(_15289_),
    .Y(_15476_));
 sky130_fd_sc_hd__and2_1 _37839_ (.A(_15471_),
    .B(_15472_),
    .X(_15477_));
 sky130_fd_sc_hd__a21o_1 _37840_ (.A1(_15456_),
    .A2(_15459_),
    .B1(_15460_),
    .X(_15478_));
 sky130_fd_sc_hd__nand3_4 _37841_ (.A(_15460_),
    .B(_15456_),
    .C(_15459_),
    .Y(_15479_));
 sky130_fd_sc_hd__nand3_2 _37842_ (.A(_15477_),
    .B(_15478_),
    .C(_15479_),
    .Y(_15480_));
 sky130_fd_sc_hd__nand3_4 _37843_ (.A(_15474_),
    .B(_15476_),
    .C(_15480_),
    .Y(_15481_));
 sky130_fd_sc_hd__o21ai_2 _37844_ (.A1(_15461_),
    .A2(_15463_),
    .B1(_15477_),
    .Y(_15482_));
 sky130_fd_sc_hd__o211a_1 _37845_ (.A1(_15024_),
    .A2(_15030_),
    .B1(_15284_),
    .C1(_15285_),
    .X(_15483_));
 sky130_fd_sc_hd__a21oi_4 _37846_ (.A1(_15287_),
    .A2(_15291_),
    .B1(_15483_),
    .Y(_15484_));
 sky130_fd_sc_hd__nand3_2 _37847_ (.A(_15478_),
    .B(_15479_),
    .C(_15473_),
    .Y(_15485_));
 sky130_fd_sc_hd__nand3_4 _37848_ (.A(_15482_),
    .B(_15484_),
    .C(_15485_),
    .Y(_15486_));
 sky130_fd_sc_hd__nand2_4 _37849_ (.A(_15347_),
    .B(_15346_),
    .Y(_15487_));
 sky130_fd_sc_hd__a21oi_2 _37850_ (.A1(_15481_),
    .A2(_15486_),
    .B1(_15487_),
    .Y(_15488_));
 sky130_fd_sc_hd__nand3_4 _37851_ (.A(_15481_),
    .B(_15486_),
    .C(_15487_),
    .Y(_15489_));
 sky130_vsdinv _37852_ (.A(_15489_),
    .Y(_15490_));
 sky130_fd_sc_hd__nand2_1 _37853_ (.A(_15251_),
    .B(_15228_),
    .Y(_15491_));
 sky130_fd_sc_hd__nand2_2 _37854_ (.A(_15491_),
    .B(_15232_),
    .Y(_15492_));
 sky130_fd_sc_hd__nand3_4 _37855_ (.A(_12780_),
    .B(_12401_),
    .C(_07323_),
    .Y(_15493_));
 sky130_fd_sc_hd__nand2_1 _37856_ (.A(_13737_),
    .B(_07323_),
    .Y(_15494_));
 sky130_fd_sc_hd__o21ai_4 _37857_ (.A1(_11848_),
    .A2(_13099_),
    .B1(_15494_),
    .Y(_15495_));
 sky130_fd_sc_hd__o21ai_2 _37858_ (.A1(net435),
    .A2(_15493_),
    .B1(_15495_),
    .Y(_15496_));
 sky130_fd_sc_hd__nand2_2 _37859_ (.A(_19580_),
    .B(_07055_),
    .Y(_15497_));
 sky130_fd_sc_hd__nand2_4 _37860_ (.A(_15496_),
    .B(_15497_),
    .Y(_15498_));
 sky130_fd_sc_hd__nor2_2 _37861_ (.A(net435),
    .B(_15493_),
    .Y(_15499_));
 sky130_vsdinv _37862_ (.A(_15497_),
    .Y(_15500_));
 sky130_fd_sc_hd__nand3b_4 _37863_ (.A_N(_15499_),
    .B(_15500_),
    .C(_15495_),
    .Y(_15501_));
 sky130_fd_sc_hd__o21ai_4 _37864_ (.A1(_15203_),
    .A2(_15209_),
    .B1(_15201_),
    .Y(_15502_));
 sky130_fd_sc_hd__a21oi_4 _37865_ (.A1(_15498_),
    .A2(_15501_),
    .B1(_15502_),
    .Y(_15503_));
 sky130_fd_sc_hd__and3_1 _37866_ (.A(_15498_),
    .B(_15502_),
    .C(_15501_),
    .X(_15504_));
 sky130_fd_sc_hd__nand2_1 _37867_ (.A(_19583_),
    .B(_08734_),
    .Y(_15505_));
 sky130_fd_sc_hd__nand2_2 _37868_ (.A(_10282_),
    .B(_08735_),
    .Y(_15506_));
 sky130_fd_sc_hd__nor2_2 _37869_ (.A(_15505_),
    .B(_15506_),
    .Y(_15507_));
 sky130_fd_sc_hd__nand2_1 _37870_ (.A(_15505_),
    .B(_15506_),
    .Y(_15508_));
 sky130_vsdinv _37871_ (.A(_15508_),
    .Y(_15509_));
 sky130_fd_sc_hd__nor2_1 _37872_ (.A(net468),
    .B(_10960_),
    .Y(_15510_));
 sky130_fd_sc_hd__o21bai_2 _37873_ (.A1(_15507_),
    .A2(_15509_),
    .B1_N(_15510_),
    .Y(_15511_));
 sky130_fd_sc_hd__nand3b_2 _37874_ (.A_N(_15507_),
    .B(_15510_),
    .C(_15508_),
    .Y(_15512_));
 sky130_fd_sc_hd__nand2_4 _37875_ (.A(_15511_),
    .B(_15512_),
    .Y(_15513_));
 sky130_vsdinv _37876_ (.A(_15513_),
    .Y(_15514_));
 sky130_fd_sc_hd__o21ai_4 _37877_ (.A1(_15503_),
    .A2(_15504_),
    .B1(_15514_),
    .Y(_15515_));
 sky130_fd_sc_hd__a21boi_4 _37878_ (.A1(_15213_),
    .A2(_15226_),
    .B1_N(_15207_),
    .Y(_15516_));
 sky130_fd_sc_hd__a21o_1 _37879_ (.A1(_15498_),
    .A2(_15501_),
    .B1(_15502_),
    .X(_15517_));
 sky130_fd_sc_hd__nand3_4 _37880_ (.A(_15498_),
    .B(_15502_),
    .C(_15501_),
    .Y(_15518_));
 sky130_fd_sc_hd__nand3_4 _37881_ (.A(_15517_),
    .B(_15518_),
    .C(_15513_),
    .Y(_15519_));
 sky130_fd_sc_hd__nand3_4 _37882_ (.A(_15515_),
    .B(_15516_),
    .C(_15519_),
    .Y(_15520_));
 sky130_fd_sc_hd__o21ai_2 _37883_ (.A1(_15503_),
    .A2(_15504_),
    .B1(_15513_),
    .Y(_15521_));
 sky130_fd_sc_hd__nand2_1 _37884_ (.A(_15213_),
    .B(_15226_),
    .Y(_15522_));
 sky130_fd_sc_hd__nand2_1 _37885_ (.A(_15522_),
    .B(_15207_),
    .Y(_15523_));
 sky130_fd_sc_hd__nand3_2 _37886_ (.A(_15514_),
    .B(_15517_),
    .C(_15518_),
    .Y(_15524_));
 sky130_fd_sc_hd__nand3_4 _37887_ (.A(_15521_),
    .B(_15523_),
    .C(_15524_),
    .Y(_15525_));
 sky130_fd_sc_hd__nand2_2 _37888_ (.A(_13514_),
    .B(_19869_),
    .Y(_15526_));
 sky130_fd_sc_hd__nand2_1 _37889_ (.A(_11379_),
    .B(_10738_),
    .Y(_15527_));
 sky130_fd_sc_hd__nor2_2 _37890_ (.A(_15526_),
    .B(_15527_),
    .Y(_15528_));
 sky130_fd_sc_hd__nor2_2 _37891_ (.A(_08580_),
    .B(_12078_),
    .Y(_15529_));
 sky130_fd_sc_hd__nand2_1 _37892_ (.A(_15526_),
    .B(_15527_),
    .Y(_15530_));
 sky130_fd_sc_hd__nand3b_4 _37893_ (.A_N(_15528_),
    .B(_15529_),
    .C(_15530_),
    .Y(_15531_));
 sky130_fd_sc_hd__a21o_1 _37894_ (.A1(_19601_),
    .A2(_10745_),
    .B1(_15526_),
    .X(_15532_));
 sky130_fd_sc_hd__a21o_1 _37895_ (.A1(_19598_),
    .A2(_11724_),
    .B1(_15527_),
    .X(_15533_));
 sky130_fd_sc_hd__o211ai_4 _37896_ (.A1(_08580_),
    .A2(_12078_),
    .B1(_15532_),
    .C1(_15533_),
    .Y(_15534_));
 sky130_fd_sc_hd__nand2_1 _37897_ (.A(_15214_),
    .B(_15215_),
    .Y(_15535_));
 sky130_fd_sc_hd__a21o_1 _37898_ (.A1(_15219_),
    .A2(_15535_),
    .B1(_15216_),
    .X(_15536_));
 sky130_fd_sc_hd__a21o_2 _37899_ (.A1(_15531_),
    .A2(_15534_),
    .B1(_15536_),
    .X(_15537_));
 sky130_fd_sc_hd__nand3_4 _37900_ (.A(_15531_),
    .B(_15536_),
    .C(_15534_),
    .Y(_15538_));
 sky130_fd_sc_hd__nand2_4 _37901_ (.A(_15244_),
    .B(_15242_),
    .Y(_15539_));
 sky130_fd_sc_hd__a21oi_4 _37902_ (.A1(_15537_),
    .A2(_15538_),
    .B1(_15539_),
    .Y(_15540_));
 sky130_fd_sc_hd__nand3_2 _37903_ (.A(_15537_),
    .B(_15539_),
    .C(_15538_),
    .Y(_15541_));
 sky130_vsdinv _37904_ (.A(_15541_),
    .Y(_15542_));
 sky130_fd_sc_hd__o2bb2ai_4 _37905_ (.A1_N(_15520_),
    .A2_N(_15525_),
    .B1(_15540_),
    .B2(_15542_),
    .Y(_15543_));
 sky130_fd_sc_hd__a21oi_2 _37906_ (.A1(_15531_),
    .A2(_15534_),
    .B1(_15536_),
    .Y(_15544_));
 sky130_fd_sc_hd__and2_1 _37907_ (.A(_15244_),
    .B(_15242_),
    .X(_15545_));
 sky130_fd_sc_hd__nor2_2 _37908_ (.A(_15544_),
    .B(_15545_),
    .Y(_15546_));
 sky130_fd_sc_hd__a21oi_4 _37909_ (.A1(_15546_),
    .A2(_15538_),
    .B1(_15540_),
    .Y(_15547_));
 sky130_fd_sc_hd__nand3_4 _37910_ (.A(_15525_),
    .B(_15520_),
    .C(_15547_),
    .Y(_15548_));
 sky130_fd_sc_hd__nand3_4 _37911_ (.A(_15492_),
    .B(_15543_),
    .C(_15548_),
    .Y(_15549_));
 sky130_fd_sc_hd__a21oi_1 _37912_ (.A1(_15214_),
    .A2(_15215_),
    .B1(_15218_),
    .Y(_15550_));
 sky130_fd_sc_hd__o211a_1 _37913_ (.A1(_15216_),
    .A2(_15550_),
    .B1(_15534_),
    .C1(_15531_),
    .X(_15551_));
 sky130_fd_sc_hd__o21ai_1 _37914_ (.A1(_15544_),
    .A2(_15551_),
    .B1(_15545_),
    .Y(_15552_));
 sky130_fd_sc_hd__nand2_2 _37915_ (.A(_15552_),
    .B(_15541_),
    .Y(_15553_));
 sky130_fd_sc_hd__a21o_1 _37916_ (.A1(_15525_),
    .A2(_15520_),
    .B1(_15553_),
    .X(_15554_));
 sky130_fd_sc_hd__a21boi_2 _37917_ (.A1(_15251_),
    .A2(_15228_),
    .B1_N(_15232_),
    .Y(_15555_));
 sky130_fd_sc_hd__nand3_2 _37918_ (.A(_15525_),
    .B(_15520_),
    .C(_15553_),
    .Y(_15556_));
 sky130_fd_sc_hd__nand3_4 _37919_ (.A(_15554_),
    .B(_15555_),
    .C(_15556_),
    .Y(_15557_));
 sky130_fd_sc_hd__nand2_2 _37920_ (.A(_12468_),
    .B(_10459_),
    .Y(_15558_));
 sky130_fd_sc_hd__nand2_2 _37921_ (.A(_19612_),
    .B(_10643_),
    .Y(_15559_));
 sky130_fd_sc_hd__nor2_2 _37922_ (.A(_15558_),
    .B(_15559_),
    .Y(_15560_));
 sky130_fd_sc_hd__and2_1 _37923_ (.A(_15558_),
    .B(_15559_),
    .X(_15561_));
 sky130_fd_sc_hd__nor2_4 _37924_ (.A(_07833_),
    .B(_11545_),
    .Y(_15562_));
 sky130_fd_sc_hd__o21bai_2 _37925_ (.A1(_15560_),
    .A2(_15561_),
    .B1_N(_15562_),
    .Y(_15563_));
 sky130_fd_sc_hd__nand2_2 _37926_ (.A(_15558_),
    .B(_15559_),
    .Y(_15564_));
 sky130_fd_sc_hd__nand3b_4 _37927_ (.A_N(_15560_),
    .B(_15562_),
    .C(_15564_),
    .Y(_15565_));
 sky130_fd_sc_hd__a21o_1 _37928_ (.A1(_15276_),
    .A2(_15275_),
    .B1(_15270_),
    .X(_15566_));
 sky130_fd_sc_hd__a21oi_2 _37929_ (.A1(_15563_),
    .A2(_15565_),
    .B1(_15566_),
    .Y(_15567_));
 sky130_fd_sc_hd__and3_1 _37930_ (.A(_15563_),
    .B(_15565_),
    .C(_15566_),
    .X(_15568_));
 sky130_fd_sc_hd__nand2_2 _37931_ (.A(_11847_),
    .B(_11909_),
    .Y(_15569_));
 sky130_fd_sc_hd__nand2_4 _37932_ (.A(_11849_),
    .B(_11178_),
    .Y(_15570_));
 sky130_fd_sc_hd__or2_1 _37933_ (.A(_15569_),
    .B(_15570_),
    .X(_15571_));
 sky130_fd_sc_hd__nand2_1 _37934_ (.A(_15569_),
    .B(_15570_),
    .Y(_15572_));
 sky130_fd_sc_hd__nand2_1 _37935_ (.A(_19629_),
    .B(_11583_),
    .Y(_15573_));
 sky130_fd_sc_hd__a21o_1 _37936_ (.A1(_15571_),
    .A2(_15572_),
    .B1(_15573_),
    .X(_15574_));
 sky130_fd_sc_hd__nand3_1 _37937_ (.A(_15571_),
    .B(_15573_),
    .C(_15572_),
    .Y(_15575_));
 sky130_fd_sc_hd__nand2_2 _37938_ (.A(_15574_),
    .B(_15575_),
    .Y(_15576_));
 sky130_fd_sc_hd__o21bai_4 _37939_ (.A1(_15567_),
    .A2(_15568_),
    .B1_N(_15576_),
    .Y(_15577_));
 sky130_fd_sc_hd__a21o_1 _37940_ (.A1(_15563_),
    .A2(_15565_),
    .B1(_15566_),
    .X(_15578_));
 sky130_fd_sc_hd__nand3_2 _37941_ (.A(_15563_),
    .B(_15565_),
    .C(_15566_),
    .Y(_15579_));
 sky130_fd_sc_hd__nand3_4 _37942_ (.A(_15578_),
    .B(_15576_),
    .C(_15579_),
    .Y(_15580_));
 sky130_fd_sc_hd__o21ai_4 _37943_ (.A1(_15246_),
    .A2(_15247_),
    .B1(_15245_),
    .Y(_15581_));
 sky130_fd_sc_hd__a21o_2 _37944_ (.A1(_15577_),
    .A2(_15580_),
    .B1(_15581_),
    .X(_15582_));
 sky130_fd_sc_hd__nand3_4 _37945_ (.A(_15577_),
    .B(_15581_),
    .C(_15580_),
    .Y(_15583_));
 sky130_vsdinv _37946_ (.A(_15279_),
    .Y(_15584_));
 sky130_fd_sc_hd__a21oi_4 _37947_ (.A1(_15283_),
    .A2(_15267_),
    .B1(_15584_),
    .Y(_15585_));
 sky130_vsdinv _37948_ (.A(_15585_),
    .Y(_15586_));
 sky130_fd_sc_hd__a21oi_4 _37949_ (.A1(_15582_),
    .A2(_15583_),
    .B1(_15586_),
    .Y(_15587_));
 sky130_fd_sc_hd__nand3_2 _37950_ (.A(_15582_),
    .B(_15583_),
    .C(_15586_),
    .Y(_15588_));
 sky130_vsdinv _37951_ (.A(_15588_),
    .Y(_15589_));
 sky130_fd_sc_hd__o2bb2ai_4 _37952_ (.A1_N(_15549_),
    .A2_N(_15557_),
    .B1(_15587_),
    .B2(_15589_),
    .Y(_15590_));
 sky130_fd_sc_hd__a21oi_4 _37953_ (.A1(_15577_),
    .A2(_15580_),
    .B1(_15581_),
    .Y(_15591_));
 sky130_fd_sc_hd__nor2_4 _37954_ (.A(_15585_),
    .B(_15591_),
    .Y(_15592_));
 sky130_fd_sc_hd__a21oi_2 _37955_ (.A1(_15583_),
    .A2(_15592_),
    .B1(_15587_),
    .Y(_15593_));
 sky130_fd_sc_hd__nand3_4 _37956_ (.A(_15593_),
    .B(_15557_),
    .C(_15549_),
    .Y(_15594_));
 sky130_fd_sc_hd__nand2_1 _37957_ (.A(_15295_),
    .B(_15257_),
    .Y(_15595_));
 sky130_fd_sc_hd__nand2_4 _37958_ (.A(_15595_),
    .B(_15261_),
    .Y(_15596_));
 sky130_fd_sc_hd__a21oi_4 _37959_ (.A1(_15590_),
    .A2(_15594_),
    .B1(_15596_),
    .Y(_15597_));
 sky130_fd_sc_hd__a21oi_4 _37960_ (.A1(_15252_),
    .A2(_15256_),
    .B1(_15254_),
    .Y(_15598_));
 sky130_fd_sc_hd__a21oi_1 _37961_ (.A1(_15285_),
    .A2(_15284_),
    .B1(_15288_),
    .Y(_15599_));
 sky130_fd_sc_hd__o21bai_1 _37962_ (.A1(_15599_),
    .A2(_15483_),
    .B1_N(_15291_),
    .Y(_15600_));
 sky130_fd_sc_hd__nand2_1 _37963_ (.A(_15600_),
    .B(_15475_),
    .Y(_15601_));
 sky130_fd_sc_hd__a31oi_4 _37964_ (.A1(_15254_),
    .A2(_15252_),
    .A3(_15256_),
    .B1(_15601_),
    .Y(_15602_));
 sky130_fd_sc_hd__o211a_2 _37965_ (.A1(_15598_),
    .A2(_15602_),
    .B1(_15594_),
    .C1(_15590_),
    .X(_15603_));
 sky130_fd_sc_hd__o22ai_4 _37966_ (.A1(_15488_),
    .A2(_15490_),
    .B1(_15597_),
    .B2(_15603_),
    .Y(_15604_));
 sky130_fd_sc_hd__o21ai_2 _37967_ (.A1(_15359_),
    .A2(_15299_),
    .B1(_15364_),
    .Y(_15605_));
 sky130_fd_sc_hd__nand2_1 _37968_ (.A(_15481_),
    .B(_15486_),
    .Y(_15606_));
 sky130_vsdinv _37969_ (.A(_15487_),
    .Y(_15607_));
 sky130_fd_sc_hd__nand2_1 _37970_ (.A(_15606_),
    .B(_15607_),
    .Y(_15608_));
 sky130_fd_sc_hd__nand2_4 _37971_ (.A(_15608_),
    .B(_15489_),
    .Y(_15609_));
 sky130_fd_sc_hd__nand2_1 _37972_ (.A(_15590_),
    .B(_15594_),
    .Y(_15610_));
 sky130_fd_sc_hd__nor2_2 _37973_ (.A(_15598_),
    .B(_15602_),
    .Y(_15611_));
 sky130_fd_sc_hd__nand2_2 _37974_ (.A(_15610_),
    .B(_15611_),
    .Y(_15612_));
 sky130_fd_sc_hd__nand3_4 _37975_ (.A(_15596_),
    .B(_15590_),
    .C(_15594_),
    .Y(_15613_));
 sky130_fd_sc_hd__nand3b_4 _37976_ (.A_N(_15609_),
    .B(_15612_),
    .C(_15613_),
    .Y(_15614_));
 sky130_fd_sc_hd__nand3_4 _37977_ (.A(_15604_),
    .B(_15605_),
    .C(_15614_),
    .Y(_15615_));
 sky130_fd_sc_hd__o21a_1 _37978_ (.A1(_15359_),
    .A2(_15299_),
    .B1(_15364_),
    .X(_15616_));
 sky130_fd_sc_hd__o21bai_2 _37979_ (.A1(_15597_),
    .A2(_15603_),
    .B1_N(_15609_),
    .Y(_15617_));
 sky130_fd_sc_hd__nand3_2 _37980_ (.A(_15612_),
    .B(_15613_),
    .C(_15609_),
    .Y(_15618_));
 sky130_fd_sc_hd__nand3_4 _37981_ (.A(_15616_),
    .B(_15617_),
    .C(_15618_),
    .Y(_15619_));
 sky130_vsdinv _37982_ (.A(_15394_),
    .Y(_15620_));
 sky130_fd_sc_hd__and2_1 _37983_ (.A(_15389_),
    .B(_13663_),
    .X(_15621_));
 sky130_fd_sc_hd__and3_1 _37984_ (.A(_15333_),
    .B(_15336_),
    .C(_15337_),
    .X(_15622_));
 sky130_fd_sc_hd__o21ai_2 _37985_ (.A1(_14815_),
    .A2(_15622_),
    .B1(_15339_),
    .Y(_15623_));
 sky130_fd_sc_hd__nand3_4 _37986_ (.A(_15623_),
    .B(_15114_),
    .C(_15113_),
    .Y(_15624_));
 sky130_fd_sc_hd__nand3_4 _37987_ (.A(_15115_),
    .B(_15339_),
    .C(_15341_),
    .Y(_15625_));
 sky130_fd_sc_hd__nand2_2 _37988_ (.A(_15624_),
    .B(_15625_),
    .Y(_15626_));
 sky130_fd_sc_hd__nand2_2 _37989_ (.A(_15626_),
    .B(_15392_),
    .Y(_15627_));
 sky130_fd_sc_hd__nand3_4 _37990_ (.A(_15624_),
    .B(_15625_),
    .C(_15381_),
    .Y(_15628_));
 sky130_fd_sc_hd__nand2_2 _37991_ (.A(_15390_),
    .B(_15379_),
    .Y(_15629_));
 sky130_fd_sc_hd__a21oi_4 _37992_ (.A1(_15627_),
    .A2(_15628_),
    .B1(_15629_),
    .Y(_15630_));
 sky130_fd_sc_hd__nand3_2 _37993_ (.A(_15627_),
    .B(_15629_),
    .C(_15628_),
    .Y(_15631_));
 sky130_vsdinv _37994_ (.A(_15631_),
    .Y(_15632_));
 sky130_fd_sc_hd__o21ai_1 _37995_ (.A1(_15630_),
    .A2(_15632_),
    .B1(_14283_),
    .Y(_15633_));
 sky130_fd_sc_hd__o21ai_1 _37996_ (.A1(_15352_),
    .A2(_15349_),
    .B1(_15357_),
    .Y(_15634_));
 sky130_fd_sc_hd__a21o_1 _37997_ (.A1(_15627_),
    .A2(_15628_),
    .B1(_15629_),
    .X(_15635_));
 sky130_fd_sc_hd__nand3_1 _37998_ (.A(_15635_),
    .B(_13988_),
    .C(_15631_),
    .Y(_15636_));
 sky130_fd_sc_hd__nand3_1 _37999_ (.A(_15633_),
    .B(_15634_),
    .C(_15636_),
    .Y(_15637_));
 sky130_fd_sc_hd__o21ai_2 _38000_ (.A1(_15630_),
    .A2(_15632_),
    .B1(_13979_),
    .Y(_15638_));
 sky130_fd_sc_hd__a21oi_4 _38001_ (.A1(_15356_),
    .A2(_15351_),
    .B1(_15350_),
    .Y(_15639_));
 sky130_fd_sc_hd__nand3_2 _38002_ (.A(_15635_),
    .B(_13656_),
    .C(_15631_),
    .Y(_15640_));
 sky130_fd_sc_hd__nand3_4 _38003_ (.A(_15638_),
    .B(_15639_),
    .C(_15640_),
    .Y(_15641_));
 sky130_fd_sc_hd__o211a_1 _38004_ (.A1(_15620_),
    .A2(_15621_),
    .B1(_15637_),
    .C1(_15641_),
    .X(_15642_));
 sky130_fd_sc_hd__clkbuf_2 _38005_ (.A(_15637_),
    .X(_15643_));
 sky130_fd_sc_hd__or2_2 _38006_ (.A(_15620_),
    .B(_15621_),
    .X(_15644_));
 sky130_fd_sc_hd__a21oi_2 _38007_ (.A1(_15641_),
    .A2(_15643_),
    .B1(_15644_),
    .Y(_15645_));
 sky130_fd_sc_hd__o2bb2ai_1 _38008_ (.A1_N(_15615_),
    .A2_N(_15619_),
    .B1(_15642_),
    .B2(_15645_),
    .Y(_15646_));
 sky130_vsdinv _38009_ (.A(_15372_),
    .Y(_15647_));
 sky130_fd_sc_hd__nand2_1 _38010_ (.A(_15370_),
    .B(_15373_),
    .Y(_15648_));
 sky130_fd_sc_hd__o2bb2ai_2 _38011_ (.A1_N(_15366_),
    .A2_N(_15409_),
    .B1(_15647_),
    .B2(_15648_),
    .Y(_15649_));
 sky130_fd_sc_hd__nor2_2 _38012_ (.A(_15645_),
    .B(_15642_),
    .Y(_15650_));
 sky130_fd_sc_hd__nand3_2 _38013_ (.A(_15650_),
    .B(_15619_),
    .C(_15615_),
    .Y(_15651_));
 sky130_fd_sc_hd__nand3_4 _38014_ (.A(_15646_),
    .B(_15649_),
    .C(_15651_),
    .Y(_15652_));
 sky130_fd_sc_hd__nand2_1 _38015_ (.A(_15619_),
    .B(_15615_),
    .Y(_15653_));
 sky130_fd_sc_hd__nand2_1 _38016_ (.A(_15653_),
    .B(_15650_),
    .Y(_15654_));
 sky130_fd_sc_hd__a21boi_4 _38017_ (.A1(_15409_),
    .A2(_15366_),
    .B1_N(_15374_),
    .Y(_15655_));
 sky130_fd_sc_hd__a21o_1 _38018_ (.A1(_15641_),
    .A2(_15643_),
    .B1(_15644_),
    .X(_15656_));
 sky130_fd_sc_hd__nand3_1 _38019_ (.A(_15644_),
    .B(_15641_),
    .C(_15643_),
    .Y(_15657_));
 sky130_fd_sc_hd__nand2_2 _38020_ (.A(_15656_),
    .B(_15657_),
    .Y(_15658_));
 sky130_fd_sc_hd__nand3_2 _38021_ (.A(_15658_),
    .B(_15619_),
    .C(_15615_),
    .Y(_15659_));
 sky130_fd_sc_hd__nand3_4 _38022_ (.A(_15654_),
    .B(_15655_),
    .C(_15659_),
    .Y(_15660_));
 sky130_fd_sc_hd__nand3_1 _38023_ (.A(_15400_),
    .B(_15403_),
    .C(_15405_),
    .Y(_15661_));
 sky130_fd_sc_hd__nand2_2 _38024_ (.A(_15661_),
    .B(_15403_),
    .Y(_15662_));
 sky130_vsdinv _38025_ (.A(_15662_),
    .Y(_15663_));
 sky130_fd_sc_hd__nor2_2 _38026_ (.A(_14595_),
    .B(_15663_),
    .Y(_15664_));
 sky130_fd_sc_hd__clkbuf_2 _38027_ (.A(_15664_),
    .X(_15665_));
 sky130_fd_sc_hd__nor2_2 _38028_ (.A(_14305_),
    .B(_15662_),
    .Y(_15666_));
 sky130_fd_sc_hd__o2bb2ai_1 _38029_ (.A1_N(_15652_),
    .A2_N(_15660_),
    .B1(_15665_),
    .B2(_15666_),
    .Y(_15667_));
 sky130_fd_sc_hd__nand2_1 _38030_ (.A(_15413_),
    .B(_15197_),
    .Y(_15668_));
 sky130_fd_sc_hd__nand2_1 _38031_ (.A(_15668_),
    .B(_15419_),
    .Y(_15669_));
 sky130_fd_sc_hd__nor2_4 _38032_ (.A(_15666_),
    .B(_15664_),
    .Y(_15670_));
 sky130_fd_sc_hd__nand3_2 _38033_ (.A(_15660_),
    .B(_15652_),
    .C(_15670_),
    .Y(_15671_));
 sky130_fd_sc_hd__nand3_4 _38034_ (.A(_15667_),
    .B(_15669_),
    .C(_15671_),
    .Y(_15672_));
 sky130_fd_sc_hd__nor2_1 _38035_ (.A(_14903_),
    .B(_15663_),
    .Y(_15673_));
 sky130_fd_sc_hd__nor2_1 _38036_ (.A(_14330_),
    .B(_15662_),
    .Y(_15674_));
 sky130_fd_sc_hd__o2bb2ai_1 _38037_ (.A1_N(_15652_),
    .A2_N(_15660_),
    .B1(_15673_),
    .B2(_15674_),
    .Y(_15675_));
 sky130_fd_sc_hd__a21boi_2 _38038_ (.A1(_15413_),
    .A2(_15197_),
    .B1_N(_15419_),
    .Y(_15676_));
 sky130_fd_sc_hd__nand3b_1 _38039_ (.A_N(_15670_),
    .B(_15660_),
    .C(_15652_),
    .Y(_15677_));
 sky130_fd_sc_hd__nand3_2 _38040_ (.A(_15675_),
    .B(_15676_),
    .C(_15677_),
    .Y(_15678_));
 sky130_fd_sc_hd__and3_2 _38041_ (.A(_15672_),
    .B(_15678_),
    .C(_15196_),
    .X(_15679_));
 sky130_fd_sc_hd__nand2_1 _38042_ (.A(_15672_),
    .B(_15678_),
    .Y(_15680_));
 sky130_vsdinv _38043_ (.A(_15196_),
    .Y(_15681_));
 sky130_fd_sc_hd__nand2_1 _38044_ (.A(_15680_),
    .B(_15681_),
    .Y(_15682_));
 sky130_fd_sc_hd__a21oi_1 _38045_ (.A1(_15426_),
    .A2(_15427_),
    .B1(_15425_),
    .Y(_15683_));
 sky130_fd_sc_hd__o21ai_2 _38046_ (.A1(_15431_),
    .A2(_15683_),
    .B1(_15428_),
    .Y(_15684_));
 sky130_fd_sc_hd__nand2_2 _38047_ (.A(_15682_),
    .B(_15684_),
    .Y(_15685_));
 sky130_fd_sc_hd__a21oi_1 _38048_ (.A1(_15672_),
    .A2(_15678_),
    .B1(_15196_),
    .Y(_15686_));
 sky130_fd_sc_hd__o21bai_2 _38049_ (.A1(_15686_),
    .A2(_15679_),
    .B1_N(_15684_),
    .Y(_15687_));
 sky130_fd_sc_hd__o21a_1 _38050_ (.A1(_15679_),
    .A2(_15685_),
    .B1(_15687_),
    .X(_15688_));
 sky130_vsdinv _38051_ (.A(_15688_),
    .Y(_15689_));
 sky130_fd_sc_hd__and4_2 _38052_ (.A(_15178_),
    .B(_15183_),
    .C(_15433_),
    .D(_15437_),
    .X(_15690_));
 sky130_fd_sc_hd__nand2_1 _38053_ (.A(_15183_),
    .B(_15437_),
    .Y(_15691_));
 sky130_fd_sc_hd__nand2_2 _38054_ (.A(_15691_),
    .B(_15433_),
    .Y(_15692_));
 sky130_fd_sc_hd__a21boi_4 _38055_ (.A1(_15190_),
    .A2(_15690_),
    .B1_N(_15692_),
    .Y(_15693_));
 sky130_fd_sc_hd__xor2_4 _38056_ (.A(_15689_),
    .B(_15693_),
    .X(_02665_));
 sky130_fd_sc_hd__nor2_1 _38057_ (.A(_15679_),
    .B(_15685_),
    .Y(_15694_));
 sky130_vsdinv _38058_ (.A(_15694_),
    .Y(_15695_));
 sky130_fd_sc_hd__o21ai_1 _38059_ (.A1(_15689_),
    .A2(_15693_),
    .B1(_15695_),
    .Y(_15696_));
 sky130_fd_sc_hd__and2_4 _38060_ (.A(_15465_),
    .B(net478),
    .X(_15697_));
 sky130_fd_sc_hd__a21oi_2 _38061_ (.A1(_15470_),
    .A2(_14809_),
    .B1(_15697_),
    .Y(_15698_));
 sky130_fd_sc_hd__nor2_4 _38062_ (.A(_13945_),
    .B(_15109_),
    .Y(_15699_));
 sky130_fd_sc_hd__nor2_4 _38063_ (.A(_14257_),
    .B(_15111_),
    .Y(_15700_));
 sky130_fd_sc_hd__nor2_1 _38064_ (.A(_15699_),
    .B(_15700_),
    .Y(_15701_));
 sky130_fd_sc_hd__nand2_2 _38065_ (.A(_15698_),
    .B(_15701_),
    .Y(_15702_));
 sky130_vsdinv _38066_ (.A(_15700_),
    .Y(_15703_));
 sky130_vsdinv _38067_ (.A(_15699_),
    .Y(_15704_));
 sky130_vsdinv _38068_ (.A(_15697_),
    .Y(_15705_));
 sky130_fd_sc_hd__a22o_1 _38069_ (.A1(_15703_),
    .A2(_15704_),
    .B1(_15471_),
    .B2(_15705_),
    .X(_15706_));
 sky130_fd_sc_hd__o2111ai_4 _38070_ (.A1(_15392_),
    .A2(_15626_),
    .B1(_15624_),
    .C1(_15702_),
    .D1(_15706_),
    .Y(_15707_));
 sky130_fd_sc_hd__nand2_1 _38071_ (.A(_15706_),
    .B(_15702_),
    .Y(_15708_));
 sky130_fd_sc_hd__nand2_1 _38072_ (.A(_15628_),
    .B(_15624_),
    .Y(_15709_));
 sky130_fd_sc_hd__nand2_2 _38073_ (.A(_15708_),
    .B(_15709_),
    .Y(_15710_));
 sky130_fd_sc_hd__a21o_1 _38074_ (.A1(_15707_),
    .A2(_15710_),
    .B1(_13988_),
    .X(_15711_));
 sky130_fd_sc_hd__nand3_4 _38075_ (.A(_15707_),
    .B(_15710_),
    .C(_13988_),
    .Y(_15712_));
 sky130_fd_sc_hd__nand2_2 _38076_ (.A(_15711_),
    .B(_15712_),
    .Y(_15713_));
 sky130_fd_sc_hd__a21boi_4 _38077_ (.A1(_15486_),
    .A2(_15487_),
    .B1_N(_15481_),
    .Y(_15714_));
 sky130_fd_sc_hd__nand2_4 _38078_ (.A(_15713_),
    .B(_15714_),
    .Y(_15715_));
 sky130_fd_sc_hd__nor2_1 _38079_ (.A(_14283_),
    .B(_15630_),
    .Y(_15716_));
 sky130_fd_sc_hd__nor2_2 _38080_ (.A(_15632_),
    .B(_15716_),
    .Y(_15717_));
 sky130_vsdinv _38081_ (.A(_15717_),
    .Y(_15718_));
 sky130_fd_sc_hd__nand2_1 _38082_ (.A(_15489_),
    .B(_15481_),
    .Y(_15719_));
 sky130_fd_sc_hd__nand3_4 _38083_ (.A(_15719_),
    .B(_15712_),
    .C(_15711_),
    .Y(_15720_));
 sky130_fd_sc_hd__nand3_1 _38084_ (.A(_15715_),
    .B(_15718_),
    .C(_15720_),
    .Y(_15721_));
 sky130_vsdinv _38085_ (.A(_15721_),
    .Y(_15722_));
 sky130_fd_sc_hd__a21oi_4 _38086_ (.A1(_15715_),
    .A2(_15720_),
    .B1(_15718_),
    .Y(_15723_));
 sky130_fd_sc_hd__and3_2 _38087_ (.A(_15577_),
    .B(_15581_),
    .C(_15580_),
    .X(_15724_));
 sky130_fd_sc_hd__nand2_1 _38088_ (.A(_19633_),
    .B(_19830_),
    .Y(_15725_));
 sky130_fd_sc_hd__nand2_2 _38089_ (.A(_10991_),
    .B(_11200_),
    .Y(_15726_));
 sky130_fd_sc_hd__nor2_1 _38090_ (.A(_15725_),
    .B(_15726_),
    .Y(_15727_));
 sky130_fd_sc_hd__and2_1 _38091_ (.A(_15725_),
    .B(_15726_),
    .X(_15728_));
 sky130_fd_sc_hd__nor2_8 _38092_ (.A(_18468_),
    .B(_06433_),
    .Y(_15729_));
 sky130_vsdinv _38093_ (.A(_15729_),
    .Y(_15730_));
 sky130_fd_sc_hd__o21ai_2 _38094_ (.A1(_15727_),
    .A2(_15728_),
    .B1(_15730_),
    .Y(_15731_));
 sky130_fd_sc_hd__or2_2 _38095_ (.A(_15725_),
    .B(_15726_),
    .X(_15732_));
 sky130_fd_sc_hd__nand2_1 _38096_ (.A(_15725_),
    .B(_15726_),
    .Y(_15733_));
 sky130_fd_sc_hd__nand3_4 _38097_ (.A(_15732_),
    .B(_15729_),
    .C(_15733_),
    .Y(_15734_));
 sky130_fd_sc_hd__nor2_1 _38098_ (.A(_15569_),
    .B(_15570_),
    .Y(_15735_));
 sky130_fd_sc_hd__a31oi_2 _38099_ (.A1(_15572_),
    .A2(_19629_),
    .A3(_19841_),
    .B1(_15735_),
    .Y(_15736_));
 sky130_fd_sc_hd__a21bo_1 _38100_ (.A1(_15731_),
    .A2(_15734_),
    .B1_N(_15736_),
    .X(_15737_));
 sky130_fd_sc_hd__nand3b_4 _38101_ (.A_N(_15736_),
    .B(_15731_),
    .C(_15734_),
    .Y(_15738_));
 sky130_fd_sc_hd__and2_1 _38102_ (.A(_15449_),
    .B(_15447_),
    .X(_15739_));
 sky130_fd_sc_hd__a21bo_2 _38103_ (.A1(_15737_),
    .A2(_15738_),
    .B1_N(_15739_),
    .X(_15740_));
 sky130_fd_sc_hd__nand3b_4 _38104_ (.A_N(_15739_),
    .B(_15738_),
    .C(_15737_),
    .Y(_15741_));
 sky130_fd_sc_hd__nand2_4 _38105_ (.A(_15462_),
    .B(_15458_),
    .Y(_15742_));
 sky130_fd_sc_hd__a21o_1 _38106_ (.A1(_15740_),
    .A2(_15741_),
    .B1(_15742_),
    .X(_15743_));
 sky130_fd_sc_hd__nand3_4 _38107_ (.A(_15740_),
    .B(_15742_),
    .C(_15741_),
    .Y(_15744_));
 sky130_fd_sc_hd__a21o_2 _38108_ (.A1(_14946_),
    .A2(_15464_),
    .B1(_15697_),
    .X(_15745_));
 sky130_fd_sc_hd__nor2_8 _38109_ (.A(_14815_),
    .B(_15745_),
    .Y(_15746_));
 sky130_fd_sc_hd__and2_2 _38110_ (.A(_15745_),
    .B(_14814_),
    .X(_15747_));
 sky130_fd_sc_hd__nor2_8 _38111_ (.A(_15746_),
    .B(_15747_),
    .Y(_15748_));
 sky130_fd_sc_hd__nand3_2 _38112_ (.A(_15743_),
    .B(_15744_),
    .C(_15748_),
    .Y(_15749_));
 sky130_fd_sc_hd__a21oi_4 _38113_ (.A1(_15740_),
    .A2(_15741_),
    .B1(_15742_),
    .Y(_15750_));
 sky130_fd_sc_hd__nor2_1 _38114_ (.A(_15452_),
    .B(_15455_),
    .Y(_15751_));
 sky130_fd_sc_hd__o211a_1 _38115_ (.A1(_15453_),
    .A2(_15751_),
    .B1(_15741_),
    .C1(_15740_),
    .X(_15752_));
 sky130_vsdinv _38116_ (.A(_15748_),
    .Y(_15753_));
 sky130_fd_sc_hd__buf_4 _38117_ (.A(_15753_),
    .X(_15754_));
 sky130_fd_sc_hd__clkbuf_4 _38118_ (.A(_15754_),
    .X(_15755_));
 sky130_fd_sc_hd__o21ai_2 _38119_ (.A1(_15750_),
    .A2(_15752_),
    .B1(_15755_),
    .Y(_15756_));
 sky130_fd_sc_hd__o211ai_4 _38120_ (.A1(_15724_),
    .A2(_15592_),
    .B1(_15749_),
    .C1(_15756_),
    .Y(_15757_));
 sky130_fd_sc_hd__clkbuf_4 _38121_ (.A(_15748_),
    .X(_15758_));
 sky130_fd_sc_hd__o21ai_2 _38122_ (.A1(_15750_),
    .A2(_15752_),
    .B1(_15758_),
    .Y(_15759_));
 sky130_fd_sc_hd__a21oi_4 _38123_ (.A1(_15582_),
    .A2(_15586_),
    .B1(_15724_),
    .Y(_15760_));
 sky130_fd_sc_hd__nand3_4 _38124_ (.A(_15743_),
    .B(_15744_),
    .C(_15754_),
    .Y(_15761_));
 sky130_fd_sc_hd__nand3_4 _38125_ (.A(_15759_),
    .B(_15760_),
    .C(_15761_),
    .Y(_15762_));
 sky130_fd_sc_hd__o21a_1 _38126_ (.A1(_15473_),
    .A2(_15461_),
    .B1(_15479_),
    .X(_15763_));
 sky130_vsdinv _38127_ (.A(_15763_),
    .Y(_15764_));
 sky130_fd_sc_hd__and3_1 _38128_ (.A(_15757_),
    .B(_15762_),
    .C(_15764_),
    .X(_15765_));
 sky130_fd_sc_hd__a21oi_4 _38129_ (.A1(_15757_),
    .A2(_15762_),
    .B1(_15764_),
    .Y(_15766_));
 sky130_fd_sc_hd__a21oi_4 _38130_ (.A1(_15537_),
    .A2(_15539_),
    .B1(_15551_),
    .Y(_15767_));
 sky130_fd_sc_hd__buf_2 _38131_ (.A(_08155_),
    .X(_15768_));
 sky130_fd_sc_hd__clkbuf_2 _38132_ (.A(_08908_),
    .X(_15769_));
 sky130_fd_sc_hd__nand2_1 _38133_ (.A(_15769_),
    .B(_19855_),
    .Y(_15770_));
 sky130_fd_sc_hd__a21o_1 _38134_ (.A1(_15768_),
    .A2(_19852_),
    .B1(_15770_),
    .X(_15771_));
 sky130_fd_sc_hd__nand2_1 _38135_ (.A(_15768_),
    .B(_11224_),
    .Y(_15772_));
 sky130_fd_sc_hd__a21o_1 _38136_ (.A1(_15769_),
    .A2(_14501_),
    .B1(_15772_),
    .X(_15773_));
 sky130_fd_sc_hd__nand2_2 _38137_ (.A(_19618_),
    .B(_15316_),
    .Y(_15774_));
 sky130_fd_sc_hd__a21o_2 _38138_ (.A1(_15771_),
    .A2(_15773_),
    .B1(_15774_),
    .X(_15775_));
 sky130_fd_sc_hd__nand3_4 _38139_ (.A(_15771_),
    .B(_15773_),
    .C(_15774_),
    .Y(_15776_));
 sky130_fd_sc_hd__a31o_2 _38140_ (.A1(_15564_),
    .A2(_19618_),
    .A3(_19853_),
    .B1(_15560_),
    .X(_15777_));
 sky130_fd_sc_hd__a21oi_4 _38141_ (.A1(_15775_),
    .A2(_15776_),
    .B1(_15777_),
    .Y(_15778_));
 sky130_fd_sc_hd__and3_2 _38142_ (.A(_15775_),
    .B(_15777_),
    .C(_15776_),
    .X(_15779_));
 sky130_fd_sc_hd__clkbuf_4 _38143_ (.A(_11206_),
    .X(_15780_));
 sky130_fd_sc_hd__nor2_4 _38144_ (.A(net471),
    .B(_15780_),
    .Y(_15781_));
 sky130_fd_sc_hd__nand2_2 _38145_ (.A(_19623_),
    .B(_19840_),
    .Y(_15782_));
 sky130_fd_sc_hd__a22o_1 _38146_ (.A1(_19623_),
    .A2(_13248_),
    .B1(_19626_),
    .B2(_11574_),
    .X(_15783_));
 sky130_fd_sc_hd__o21ai_4 _38147_ (.A1(_15570_),
    .A2(_15782_),
    .B1(_15783_),
    .Y(_15784_));
 sky130_fd_sc_hd__xor2_4 _38148_ (.A(_15781_),
    .B(_15784_),
    .X(_15785_));
 sky130_fd_sc_hd__o21ai_2 _38149_ (.A1(_15778_),
    .A2(_15779_),
    .B1(_15785_),
    .Y(_15786_));
 sky130_fd_sc_hd__a21o_1 _38150_ (.A1(_15775_),
    .A2(_15776_),
    .B1(_15777_),
    .X(_15787_));
 sky130_fd_sc_hd__nand3_2 _38151_ (.A(_15775_),
    .B(_15777_),
    .C(_15776_),
    .Y(_15788_));
 sky130_fd_sc_hd__nand3b_2 _38152_ (.A_N(_15785_),
    .B(_15787_),
    .C(_15788_),
    .Y(_15789_));
 sky130_fd_sc_hd__nand3b_4 _38153_ (.A_N(_15767_),
    .B(_15786_),
    .C(_15789_),
    .Y(_15790_));
 sky130_fd_sc_hd__o21bai_2 _38154_ (.A1(_15778_),
    .A2(_15779_),
    .B1_N(_15785_),
    .Y(_15791_));
 sky130_fd_sc_hd__nand3_2 _38155_ (.A(_15787_),
    .B(_15788_),
    .C(_15785_),
    .Y(_15792_));
 sky130_fd_sc_hd__nand3_4 _38156_ (.A(_15791_),
    .B(_15767_),
    .C(_15792_),
    .Y(_15793_));
 sky130_fd_sc_hd__a21o_2 _38157_ (.A1(_15578_),
    .A2(_15576_),
    .B1(_15568_),
    .X(_15794_));
 sky130_fd_sc_hd__and3_2 _38158_ (.A(_15790_),
    .B(_15793_),
    .C(_15794_),
    .X(_15795_));
 sky130_fd_sc_hd__a21oi_4 _38159_ (.A1(_15790_),
    .A2(_15793_),
    .B1(_15794_),
    .Y(_15796_));
 sky130_fd_sc_hd__nand2_1 _38160_ (.A(_14087_),
    .B(_10745_),
    .Y(_15797_));
 sky130_fd_sc_hd__nand2_1 _38161_ (.A(_11379_),
    .B(_19863_),
    .Y(_15798_));
 sky130_fd_sc_hd__and2_1 _38162_ (.A(_15797_),
    .B(_15798_),
    .X(_15799_));
 sky130_fd_sc_hd__nor2_1 _38163_ (.A(_15797_),
    .B(_15798_),
    .Y(_15800_));
 sky130_vsdinv _38164_ (.A(_15800_),
    .Y(_15801_));
 sky130_fd_sc_hd__buf_2 _38165_ (.A(_10466_),
    .X(_15802_));
 sky130_fd_sc_hd__nor2_2 _38166_ (.A(_08580_),
    .B(_15802_),
    .Y(_15803_));
 sky130_fd_sc_hd__nand3b_4 _38167_ (.A_N(_15799_),
    .B(_15801_),
    .C(_15803_),
    .Y(_15804_));
 sky130_fd_sc_hd__o21bai_2 _38168_ (.A1(_15800_),
    .A2(_15799_),
    .B1_N(_15803_),
    .Y(_15805_));
 sky130_fd_sc_hd__clkbuf_4 _38169_ (.A(_19592_),
    .X(_15806_));
 sky130_fd_sc_hd__a31o_2 _38170_ (.A1(_15508_),
    .A2(_15806_),
    .A3(_19872_),
    .B1(_15507_),
    .X(_15807_));
 sky130_fd_sc_hd__a21o_1 _38171_ (.A1(_15804_),
    .A2(_15805_),
    .B1(_15807_),
    .X(_15808_));
 sky130_fd_sc_hd__nand3_4 _38172_ (.A(_15804_),
    .B(_15805_),
    .C(_15807_),
    .Y(_15809_));
 sky130_vsdinv _38173_ (.A(_15531_),
    .Y(_15810_));
 sky130_fd_sc_hd__nor2_2 _38174_ (.A(_15528_),
    .B(_15810_),
    .Y(_15811_));
 sky130_fd_sc_hd__a21boi_2 _38175_ (.A1(_15808_),
    .A2(_15809_),
    .B1_N(_15811_),
    .Y(_15812_));
 sky130_fd_sc_hd__o211a_1 _38176_ (.A1(_15528_),
    .A2(_15810_),
    .B1(_15809_),
    .C1(_15808_),
    .X(_15813_));
 sky130_fd_sc_hd__buf_4 _38177_ (.A(_10286_),
    .X(_15814_));
 sky130_fd_sc_hd__nand3_4 _38178_ (.A(_13107_),
    .B(_12779_),
    .C(_06804_),
    .Y(_15815_));
 sky130_fd_sc_hd__nor2_4 _38179_ (.A(_19885_),
    .B(_15815_),
    .Y(_15816_));
 sky130_fd_sc_hd__clkbuf_2 _38180_ (.A(_11338_),
    .X(_15817_));
 sky130_fd_sc_hd__o22a_2 _38181_ (.A1(_19885_),
    .A2(_18475_),
    .B1(_15817_),
    .B2(_10993_),
    .X(_15818_));
 sky130_fd_sc_hd__o22ai_4 _38182_ (.A1(_15814_),
    .A2(net438),
    .B1(_15816_),
    .B2(_15818_),
    .Y(_15819_));
 sky130_fd_sc_hd__a21o_1 _38183_ (.A1(_15495_),
    .A2(_15500_),
    .B1(_15499_),
    .X(_15820_));
 sky130_fd_sc_hd__clkbuf_4 _38184_ (.A(_13737_),
    .X(_15821_));
 sky130_fd_sc_hd__a22o_2 _38185_ (.A1(_15821_),
    .A2(net454),
    .B1(_08007_),
    .B2(_11293_),
    .X(_15822_));
 sky130_fd_sc_hd__buf_6 _38186_ (.A(_10286_),
    .X(_15823_));
 sky130_fd_sc_hd__nor2_4 _38187_ (.A(_15823_),
    .B(net438),
    .Y(_15824_));
 sky130_fd_sc_hd__nand3b_4 _38188_ (.A_N(_15816_),
    .B(_15822_),
    .C(_15824_),
    .Y(_15825_));
 sky130_fd_sc_hd__nand3_4 _38189_ (.A(_15819_),
    .B(_15820_),
    .C(_15825_),
    .Y(_15826_));
 sky130_fd_sc_hd__o21ai_2 _38190_ (.A1(_15816_),
    .A2(_15818_),
    .B1(_15824_),
    .Y(_15827_));
 sky130_fd_sc_hd__a21oi_2 _38191_ (.A1(_15495_),
    .A2(_15500_),
    .B1(_15499_),
    .Y(_15828_));
 sky130_fd_sc_hd__o221ai_4 _38192_ (.A1(_15814_),
    .A2(net438),
    .B1(_19885_),
    .B2(_15815_),
    .C1(_15822_),
    .Y(_15829_));
 sky130_fd_sc_hd__nand3_4 _38193_ (.A(_15827_),
    .B(_15828_),
    .C(_15829_),
    .Y(_15830_));
 sky130_fd_sc_hd__nand2_2 _38194_ (.A(_19593_),
    .B(_19870_),
    .Y(_15831_));
 sky130_fd_sc_hd__and4_4 _38195_ (.A(_19584_),
    .B(_19588_),
    .C(_19872_),
    .D(_14452_),
    .X(_15832_));
 sky130_vsdinv _38196_ (.A(_11094_),
    .Y(_15833_));
 sky130_fd_sc_hd__clkbuf_4 _38197_ (.A(_15833_),
    .X(_15834_));
 sky130_fd_sc_hd__nand2_1 _38198_ (.A(_19584_),
    .B(_14452_),
    .Y(_15835_));
 sky130_fd_sc_hd__o21a_1 _38199_ (.A1(_15834_),
    .A2(_10971_),
    .B1(_15835_),
    .X(_15836_));
 sky130_fd_sc_hd__nor3_4 _38200_ (.A(_15831_),
    .B(_15832_),
    .C(_15836_),
    .Y(_15837_));
 sky130_fd_sc_hd__o21a_1 _38201_ (.A1(_15832_),
    .A2(_15836_),
    .B1(_15831_),
    .X(_15838_));
 sky130_fd_sc_hd__o2bb2ai_4 _38202_ (.A1_N(_15826_),
    .A2_N(_15830_),
    .B1(_15837_),
    .B2(_15838_),
    .Y(_15839_));
 sky130_vsdinv _38203_ (.A(_15831_),
    .Y(_15840_));
 sky130_fd_sc_hd__o21ai_1 _38204_ (.A1(_15832_),
    .A2(_15836_),
    .B1(_15840_),
    .Y(_15841_));
 sky130_fd_sc_hd__o21ai_1 _38205_ (.A1(_15834_),
    .A2(_10971_),
    .B1(_15835_),
    .Y(_15842_));
 sky130_fd_sc_hd__nand3b_1 _38206_ (.A_N(_15832_),
    .B(_15831_),
    .C(_15842_),
    .Y(_15843_));
 sky130_fd_sc_hd__nand2_2 _38207_ (.A(_15841_),
    .B(_15843_),
    .Y(_15844_));
 sky130_fd_sc_hd__nand3_4 _38208_ (.A(_15830_),
    .B(_15826_),
    .C(_15844_),
    .Y(_15845_));
 sky130_fd_sc_hd__o21ai_4 _38209_ (.A1(_15513_),
    .A2(_15503_),
    .B1(_15518_),
    .Y(_15846_));
 sky130_fd_sc_hd__a21oi_2 _38210_ (.A1(_15839_),
    .A2(_15845_),
    .B1(_15846_),
    .Y(_15847_));
 sky130_fd_sc_hd__and3_1 _38211_ (.A(_15819_),
    .B(_15820_),
    .C(_15825_),
    .X(_15848_));
 sky130_fd_sc_hd__nand2_2 _38212_ (.A(_15830_),
    .B(_15844_),
    .Y(_15849_));
 sky130_fd_sc_hd__o211a_1 _38213_ (.A1(_15848_),
    .A2(_15849_),
    .B1(_15839_),
    .C1(_15846_),
    .X(_15850_));
 sky130_fd_sc_hd__o22ai_4 _38214_ (.A1(_15812_),
    .A2(_15813_),
    .B1(_15847_),
    .B2(_15850_),
    .Y(_15851_));
 sky130_fd_sc_hd__a21oi_2 _38215_ (.A1(_15808_),
    .A2(_15809_),
    .B1(_15811_),
    .Y(_15852_));
 sky130_fd_sc_hd__and3_1 _38216_ (.A(_15808_),
    .B(_15811_),
    .C(_15809_),
    .X(_15853_));
 sky130_fd_sc_hd__nand3_4 _38217_ (.A(_15846_),
    .B(_15839_),
    .C(_15845_),
    .Y(_15854_));
 sky130_fd_sc_hd__a21o_1 _38218_ (.A1(_15839_),
    .A2(_15845_),
    .B1(_15846_),
    .X(_15855_));
 sky130_fd_sc_hd__o211ai_4 _38219_ (.A1(_15852_),
    .A2(_15853_),
    .B1(_15854_),
    .C1(_15855_),
    .Y(_15856_));
 sky130_fd_sc_hd__nand2_1 _38220_ (.A(_15520_),
    .B(_15547_),
    .Y(_15857_));
 sky130_fd_sc_hd__nand2_4 _38221_ (.A(_15857_),
    .B(_15525_),
    .Y(_15858_));
 sky130_fd_sc_hd__a21oi_4 _38222_ (.A1(_15851_),
    .A2(_15856_),
    .B1(_15858_),
    .Y(_15859_));
 sky130_fd_sc_hd__a21oi_1 _38223_ (.A1(_15515_),
    .A2(_15519_),
    .B1(_15516_),
    .Y(_15860_));
 sky130_fd_sc_hd__a31oi_1 _38224_ (.A1(_15515_),
    .A2(_15516_),
    .A3(_15519_),
    .B1(_15553_),
    .Y(_15861_));
 sky130_fd_sc_hd__o211a_2 _38225_ (.A1(_15860_),
    .A2(_15861_),
    .B1(_15856_),
    .C1(_15851_),
    .X(_15862_));
 sky130_fd_sc_hd__o22ai_4 _38226_ (.A1(_15795_),
    .A2(_15796_),
    .B1(_15859_),
    .B2(_15862_),
    .Y(_15863_));
 sky130_fd_sc_hd__a21o_1 _38227_ (.A1(_15851_),
    .A2(_15856_),
    .B1(_15858_),
    .X(_15864_));
 sky130_fd_sc_hd__nor2_4 _38228_ (.A(_15796_),
    .B(_15795_),
    .Y(_15865_));
 sky130_fd_sc_hd__nand3_4 _38229_ (.A(_15858_),
    .B(_15851_),
    .C(_15856_),
    .Y(_15866_));
 sky130_fd_sc_hd__nand3_4 _38230_ (.A(_15864_),
    .B(_15865_),
    .C(_15866_),
    .Y(_15867_));
 sky130_fd_sc_hd__o21ai_1 _38231_ (.A1(_15591_),
    .A2(_15724_),
    .B1(_15585_),
    .Y(_15868_));
 sky130_fd_sc_hd__nand2_1 _38232_ (.A(_15868_),
    .B(_15588_),
    .Y(_15869_));
 sky130_fd_sc_hd__a21oi_4 _38233_ (.A1(_15543_),
    .A2(_15548_),
    .B1(_15492_),
    .Y(_15870_));
 sky130_fd_sc_hd__o21ai_4 _38234_ (.A1(_15869_),
    .A2(_15870_),
    .B1(_15549_),
    .Y(_15871_));
 sky130_fd_sc_hd__a21oi_2 _38235_ (.A1(_15863_),
    .A2(_15867_),
    .B1(_15871_),
    .Y(_15872_));
 sky130_fd_sc_hd__nand2_1 _38236_ (.A(_15865_),
    .B(_15866_),
    .Y(_15873_));
 sky130_fd_sc_hd__o211a_1 _38237_ (.A1(_15859_),
    .A2(_15873_),
    .B1(_15863_),
    .C1(_15871_),
    .X(_15874_));
 sky130_fd_sc_hd__o22ai_4 _38238_ (.A1(_15765_),
    .A2(_15766_),
    .B1(_15872_),
    .B2(_15874_),
    .Y(_15875_));
 sky130_fd_sc_hd__a21o_1 _38239_ (.A1(_15863_),
    .A2(_15867_),
    .B1(_15871_),
    .X(_15876_));
 sky130_fd_sc_hd__a31oi_2 _38240_ (.A1(_15759_),
    .A2(_15760_),
    .A3(_15761_),
    .B1(_15763_),
    .Y(_15877_));
 sky130_fd_sc_hd__a21oi_2 _38241_ (.A1(_15757_),
    .A2(_15877_),
    .B1(_15766_),
    .Y(_15878_));
 sky130_fd_sc_hd__nand3_4 _38242_ (.A(_15871_),
    .B(_15863_),
    .C(_15867_),
    .Y(_15879_));
 sky130_fd_sc_hd__nand3_4 _38243_ (.A(_15876_),
    .B(_15878_),
    .C(_15879_),
    .Y(_15880_));
 sky130_fd_sc_hd__o21ai_4 _38244_ (.A1(_15609_),
    .A2(_15597_),
    .B1(_15613_),
    .Y(_15881_));
 sky130_fd_sc_hd__a21oi_4 _38245_ (.A1(_15875_),
    .A2(_15880_),
    .B1(_15881_),
    .Y(_15882_));
 sky130_fd_sc_hd__a21oi_1 _38246_ (.A1(_15610_),
    .A2(_15611_),
    .B1(_15609_),
    .Y(_15883_));
 sky130_fd_sc_hd__o211a_1 _38247_ (.A1(_15603_),
    .A2(_15883_),
    .B1(_15880_),
    .C1(_15875_),
    .X(_15884_));
 sky130_fd_sc_hd__o22ai_4 _38248_ (.A1(_15722_),
    .A2(_15723_),
    .B1(_15882_),
    .B2(_15884_),
    .Y(_15885_));
 sky130_fd_sc_hd__a21oi_1 _38249_ (.A1(_15604_),
    .A2(_15614_),
    .B1(_15605_),
    .Y(_15886_));
 sky130_fd_sc_hd__o21ai_2 _38250_ (.A1(_15658_),
    .A2(_15886_),
    .B1(_15615_),
    .Y(_15887_));
 sky130_fd_sc_hd__a21o_1 _38251_ (.A1(_15875_),
    .A2(_15880_),
    .B1(_15881_),
    .X(_15888_));
 sky130_fd_sc_hd__nor2_2 _38252_ (.A(_15714_),
    .B(_15713_),
    .Y(_15889_));
 sky130_fd_sc_hd__nor2_2 _38253_ (.A(_15717_),
    .B(_15889_),
    .Y(_15890_));
 sky130_fd_sc_hd__a21oi_4 _38254_ (.A1(_15890_),
    .A2(_15715_),
    .B1(_15723_),
    .Y(_15891_));
 sky130_fd_sc_hd__nand3_4 _38255_ (.A(_15875_),
    .B(_15880_),
    .C(_15881_),
    .Y(_15892_));
 sky130_fd_sc_hd__nand3_2 _38256_ (.A(_15888_),
    .B(_15891_),
    .C(_15892_),
    .Y(_15893_));
 sky130_fd_sc_hd__nand3_4 _38257_ (.A(_15885_),
    .B(_15887_),
    .C(_15893_),
    .Y(_15894_));
 sky130_fd_sc_hd__o21ai_2 _38258_ (.A1(_15882_),
    .A2(_15884_),
    .B1(_15891_),
    .Y(_15895_));
 sky130_fd_sc_hd__a21boi_2 _38259_ (.A1(_15650_),
    .A2(_15619_),
    .B1_N(_15615_),
    .Y(_15896_));
 sky130_fd_sc_hd__o211ai_2 _38260_ (.A1(_15722_),
    .A2(_15723_),
    .B1(_15892_),
    .C1(_15888_),
    .Y(_15897_));
 sky130_fd_sc_hd__nand3_4 _38261_ (.A(_15895_),
    .B(_15896_),
    .C(_15897_),
    .Y(_15898_));
 sky130_fd_sc_hd__nand2_1 _38262_ (.A(_15644_),
    .B(_15641_),
    .Y(_15899_));
 sky130_fd_sc_hd__and2_2 _38263_ (.A(_15899_),
    .B(_15643_),
    .X(_15900_));
 sky130_fd_sc_hd__nor2_8 _38264_ (.A(net411),
    .B(_15900_),
    .Y(_15901_));
 sky130_fd_sc_hd__and3_1 _38265_ (.A(_15899_),
    .B(net411),
    .C(_15643_),
    .X(_15902_));
 sky130_fd_sc_hd__o2bb2ai_2 _38266_ (.A1_N(_15894_),
    .A2_N(_15898_),
    .B1(_15901_),
    .B2(_15902_),
    .Y(_15903_));
 sky130_fd_sc_hd__nand2_1 _38267_ (.A(_15660_),
    .B(_15670_),
    .Y(_15904_));
 sky130_fd_sc_hd__nand2_1 _38268_ (.A(_15904_),
    .B(_15652_),
    .Y(_15905_));
 sky130_fd_sc_hd__nor2_4 _38269_ (.A(_15902_),
    .B(_15901_),
    .Y(_15906_));
 sky130_fd_sc_hd__nand3_2 _38270_ (.A(_15898_),
    .B(_15894_),
    .C(_15906_),
    .Y(_15907_));
 sky130_fd_sc_hd__nand3_4 _38271_ (.A(_15903_),
    .B(_15905_),
    .C(_15907_),
    .Y(_15908_));
 sky130_fd_sc_hd__nor2_1 _38272_ (.A(_14903_),
    .B(_15900_),
    .Y(_15909_));
 sky130_fd_sc_hd__and3_1 _38273_ (.A(_15899_),
    .B(_14592_),
    .C(_15643_),
    .X(_15910_));
 sky130_fd_sc_hd__o2bb2ai_2 _38274_ (.A1_N(_15894_),
    .A2_N(_15898_),
    .B1(_15909_),
    .B2(_15910_),
    .Y(_15911_));
 sky130_fd_sc_hd__a21boi_2 _38275_ (.A1(_15660_),
    .A2(_15670_),
    .B1_N(_15652_),
    .Y(_15912_));
 sky130_fd_sc_hd__nand3b_2 _38276_ (.A_N(_15906_),
    .B(_15898_),
    .C(_15894_),
    .Y(_15913_));
 sky130_fd_sc_hd__nand3_4 _38277_ (.A(_15911_),
    .B(_15912_),
    .C(_15913_),
    .Y(_15914_));
 sky130_fd_sc_hd__a21oi_2 _38278_ (.A1(_15908_),
    .A2(_15914_),
    .B1(_15665_),
    .Y(_15915_));
 sky130_fd_sc_hd__and3_1 _38279_ (.A(_15908_),
    .B(_15914_),
    .C(_15665_),
    .X(_15916_));
 sky130_fd_sc_hd__nand2_1 _38280_ (.A(_15678_),
    .B(_15196_),
    .Y(_15917_));
 sky130_fd_sc_hd__nand2_2 _38281_ (.A(_15917_),
    .B(_15672_),
    .Y(_15918_));
 sky130_fd_sc_hd__o21bai_4 _38282_ (.A1(_15915_),
    .A2(_15916_),
    .B1_N(_15918_),
    .Y(_15919_));
 sky130_fd_sc_hd__a21o_1 _38283_ (.A1(_15908_),
    .A2(_15914_),
    .B1(_15665_),
    .X(_15920_));
 sky130_fd_sc_hd__nand3_2 _38284_ (.A(_15908_),
    .B(_15914_),
    .C(_15665_),
    .Y(_15921_));
 sky130_fd_sc_hd__nand3_4 _38285_ (.A(_15920_),
    .B(_15918_),
    .C(_15921_),
    .Y(_15922_));
 sky130_fd_sc_hd__and2_2 _38286_ (.A(_15919_),
    .B(_15922_),
    .X(_15923_));
 sky130_vsdinv _38287_ (.A(_15923_),
    .Y(_15924_));
 sky130_fd_sc_hd__nand2_1 _38288_ (.A(_15696_),
    .B(_15924_),
    .Y(_15925_));
 sky130_fd_sc_hd__o211ai_2 _38289_ (.A1(_15689_),
    .A2(_15693_),
    .B1(_15695_),
    .C1(_15923_),
    .Y(_15926_));
 sky130_fd_sc_hd__nand2_2 _38290_ (.A(_15925_),
    .B(_15926_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _38291_ (.A(_19593_),
    .B(_19867_),
    .Y(_15927_));
 sky130_fd_sc_hd__nand2_4 _38292_ (.A(net469),
    .B(_11094_),
    .Y(_15928_));
 sky130_vsdinv _38293_ (.A(_15928_),
    .Y(_15929_));
 sky130_fd_sc_hd__clkbuf_2 _38294_ (.A(_15929_),
    .X(_15930_));
 sky130_vsdinv _38295_ (.A(net469),
    .Y(_15931_));
 sky130_fd_sc_hd__clkbuf_2 _38296_ (.A(_15833_),
    .X(_15932_));
 sky130_fd_sc_hd__o22a_1 _38297_ (.A1(_15931_),
    .A2(_10960_),
    .B1(_15932_),
    .B2(_10654_),
    .X(_15933_));
 sky130_fd_sc_hd__a31o_1 _38298_ (.A1(_19870_),
    .A2(_19872_),
    .A3(_15930_),
    .B1(_15933_),
    .X(_15934_));
 sky130_fd_sc_hd__nor2_1 _38299_ (.A(_15927_),
    .B(_15934_),
    .Y(_15935_));
 sky130_fd_sc_hd__and2_1 _38300_ (.A(_15934_),
    .B(_15927_),
    .X(_15936_));
 sky130_fd_sc_hd__clkbuf_2 _38301_ (.A(_12402_),
    .X(_15937_));
 sky130_fd_sc_hd__and4_2 _38302_ (.A(_10993_),
    .B(_15937_),
    .C(_15821_),
    .D(_19879_),
    .X(_15938_));
 sky130_fd_sc_hd__buf_2 _38303_ (.A(_11338_),
    .X(_15939_));
 sky130_fd_sc_hd__o22a_2 _38304_ (.A1(net454),
    .A2(_18475_),
    .B1(_15939_),
    .B2(net438),
    .X(_15940_));
 sky130_fd_sc_hd__nor2_2 _38305_ (.A(_15938_),
    .B(_15940_),
    .Y(_15941_));
 sky130_fd_sc_hd__nand3_4 _38306_ (.A(_15941_),
    .B(_19581_),
    .C(_19875_),
    .Y(_15942_));
 sky130_fd_sc_hd__nand2_1 _38307_ (.A(_19580_),
    .B(_19875_),
    .Y(_15943_));
 sky130_fd_sc_hd__o21ai_2 _38308_ (.A1(_15938_),
    .A2(_15940_),
    .B1(_15943_),
    .Y(_15944_));
 sky130_fd_sc_hd__a21o_1 _38309_ (.A1(_15822_),
    .A2(_15824_),
    .B1(_15816_),
    .X(_15945_));
 sky130_fd_sc_hd__nand3_4 _38310_ (.A(_15942_),
    .B(_15944_),
    .C(_15945_),
    .Y(_15946_));
 sky130_fd_sc_hd__a21o_1 _38311_ (.A1(_15942_),
    .A2(_15944_),
    .B1(_15945_),
    .X(_15947_));
 sky130_fd_sc_hd__a2bb2o_2 _38312_ (.A1_N(_15935_),
    .A2_N(_15936_),
    .B1(_15946_),
    .B2(_15947_),
    .X(_15948_));
 sky130_fd_sc_hd__nor2_2 _38313_ (.A(_15935_),
    .B(_15936_),
    .Y(_15949_));
 sky130_fd_sc_hd__nand3_4 _38314_ (.A(_15949_),
    .B(_15947_),
    .C(_15946_),
    .Y(_15950_));
 sky130_fd_sc_hd__nand2_4 _38315_ (.A(_15849_),
    .B(_15826_),
    .Y(_15951_));
 sky130_fd_sc_hd__a21oi_4 _38316_ (.A1(_15948_),
    .A2(_15950_),
    .B1(_15951_),
    .Y(_15952_));
 sky130_fd_sc_hd__and3_1 _38317_ (.A(_15948_),
    .B(_15951_),
    .C(_15950_),
    .X(_15953_));
 sky130_fd_sc_hd__nand2_1 _38318_ (.A(_19604_),
    .B(_19856_),
    .Y(_15954_));
 sky130_fd_sc_hd__and4_2 _38319_ (.A(_14087_),
    .B(_14084_),
    .C(_13413_),
    .D(_10981_),
    .X(_15955_));
 sky130_vsdinv _38320_ (.A(_09485_),
    .Y(_15956_));
 sky130_vsdinv _38321_ (.A(_09723_),
    .Y(_15957_));
 sky130_fd_sc_hd__o22a_1 _38322_ (.A1(_15956_),
    .A2(net439),
    .B1(_15957_),
    .B2(_15802_),
    .X(_15958_));
 sky130_fd_sc_hd__or3_4 _38323_ (.A(_15954_),
    .B(_15955_),
    .C(_15958_),
    .X(_15959_));
 sky130_fd_sc_hd__o21ai_2 _38324_ (.A1(_15955_),
    .A2(_15958_),
    .B1(_15954_),
    .Y(_15960_));
 sky130_fd_sc_hd__nand2_2 _38325_ (.A(_15959_),
    .B(_15960_),
    .Y(_15961_));
 sky130_fd_sc_hd__nor2_8 _38326_ (.A(_15832_),
    .B(_15837_),
    .Y(_15962_));
 sky130_fd_sc_hd__nand2_4 _38327_ (.A(_15961_),
    .B(_15962_),
    .Y(_15963_));
 sky130_fd_sc_hd__nand3b_4 _38328_ (.A_N(_15962_),
    .B(_15960_),
    .C(_15959_),
    .Y(_15964_));
 sky130_fd_sc_hd__nand2_4 _38329_ (.A(_15804_),
    .B(_15801_),
    .Y(_15965_));
 sky130_fd_sc_hd__a21oi_4 _38330_ (.A1(_15963_),
    .A2(_15964_),
    .B1(_15965_),
    .Y(_15966_));
 sky130_fd_sc_hd__and3_2 _38331_ (.A(_15963_),
    .B(_15965_),
    .C(_15964_),
    .X(_15967_));
 sky130_fd_sc_hd__nor2_4 _38332_ (.A(_15966_),
    .B(_15967_),
    .Y(_15968_));
 sky130_fd_sc_hd__o21ai_2 _38333_ (.A1(_15952_),
    .A2(_15953_),
    .B1(_15968_),
    .Y(_15969_));
 sky130_fd_sc_hd__nand2_2 _38334_ (.A(_15856_),
    .B(_15854_),
    .Y(_15970_));
 sky130_vsdinv _38335_ (.A(_15970_),
    .Y(_15971_));
 sky130_fd_sc_hd__a21o_1 _38336_ (.A1(_15948_),
    .A2(_15950_),
    .B1(_15951_),
    .X(_15972_));
 sky130_fd_sc_hd__nand3_4 _38337_ (.A(_15948_),
    .B(_15951_),
    .C(_15950_),
    .Y(_15973_));
 sky130_fd_sc_hd__and2_1 _38338_ (.A(_15964_),
    .B(_15965_),
    .X(_15974_));
 sky130_fd_sc_hd__a21o_1 _38339_ (.A1(_15974_),
    .A2(_15963_),
    .B1(_15966_),
    .X(_15975_));
 sky130_fd_sc_hd__nand3_2 _38340_ (.A(_15972_),
    .B(_15973_),
    .C(_15975_),
    .Y(_15976_));
 sky130_fd_sc_hd__nand3_4 _38341_ (.A(_15969_),
    .B(_15971_),
    .C(_15976_),
    .Y(_15977_));
 sky130_fd_sc_hd__o22ai_4 _38342_ (.A1(_15967_),
    .A2(_15966_),
    .B1(_15952_),
    .B2(_15953_),
    .Y(_15978_));
 sky130_fd_sc_hd__nand3_4 _38343_ (.A(_15972_),
    .B(_15973_),
    .C(_15968_),
    .Y(_15979_));
 sky130_fd_sc_hd__nand3_4 _38344_ (.A(_15978_),
    .B(_15970_),
    .C(_15979_),
    .Y(_15980_));
 sky130_fd_sc_hd__nand2_1 _38345_ (.A(_15977_),
    .B(_15980_),
    .Y(_15981_));
 sky130_fd_sc_hd__and4_1 _38346_ (.A(_19609_),
    .B(_19613_),
    .C(_15316_),
    .D(_19852_),
    .X(_15982_));
 sky130_fd_sc_hd__nand2_1 _38347_ (.A(_19619_),
    .B(_19845_),
    .Y(_15983_));
 sky130_fd_sc_hd__a22o_1 _38348_ (.A1(_19609_),
    .A2(_19853_),
    .B1(_19613_),
    .B2(_19850_),
    .X(_15984_));
 sky130_fd_sc_hd__or3b_4 _38349_ (.A(_15982_),
    .B(_15983_),
    .C_N(_15984_),
    .X(_15985_));
 sky130_vsdinv _38350_ (.A(_15984_),
    .Y(_15986_));
 sky130_fd_sc_hd__o21ai_2 _38351_ (.A1(_15982_),
    .A2(_15986_),
    .B1(_15983_),
    .Y(_15987_));
 sky130_fd_sc_hd__o21ai_2 _38352_ (.A1(_15770_),
    .A2(_15772_),
    .B1(_15775_),
    .Y(_15988_));
 sky130_fd_sc_hd__a21o_1 _38353_ (.A1(_15985_),
    .A2(_15987_),
    .B1(_15988_),
    .X(_15989_));
 sky130_fd_sc_hd__nand3_4 _38354_ (.A(_15985_),
    .B(_15987_),
    .C(_15988_),
    .Y(_15990_));
 sky130_fd_sc_hd__nand2_4 _38355_ (.A(_19629_),
    .B(_19831_),
    .Y(_15991_));
 sky130_vsdinv _38356_ (.A(_19623_),
    .Y(_15992_));
 sky130_vsdinv _38357_ (.A(_08567_),
    .Y(_15993_));
 sky130_fd_sc_hd__nor2_1 _38358_ (.A(_15992_),
    .B(_15993_),
    .Y(_15994_));
 sky130_fd_sc_hd__nand2_2 _38359_ (.A(_19626_),
    .B(_11582_),
    .Y(_15995_));
 sky130_fd_sc_hd__a32o_4 _38360_ (.A1(_15994_),
    .A2(_11582_),
    .A3(_19841_),
    .B1(_15782_),
    .B2(_15995_),
    .X(_15996_));
 sky130_fd_sc_hd__xor2_4 _38361_ (.A(_15991_),
    .B(_15996_),
    .X(_15997_));
 sky130_fd_sc_hd__a21o_2 _38362_ (.A1(_15989_),
    .A2(_15990_),
    .B1(_15997_),
    .X(_15998_));
 sky130_fd_sc_hd__nand3_4 _38363_ (.A(_15989_),
    .B(_15997_),
    .C(_15990_),
    .Y(_15999_));
 sky130_fd_sc_hd__nand2_1 _38364_ (.A(_15811_),
    .B(_15809_),
    .Y(_16000_));
 sky130_fd_sc_hd__and2_2 _38365_ (.A(_16000_),
    .B(_15808_),
    .X(_16001_));
 sky130_fd_sc_hd__a21o_1 _38366_ (.A1(_15998_),
    .A2(_15999_),
    .B1(_16001_),
    .X(_16002_));
 sky130_fd_sc_hd__nand3_4 _38367_ (.A(_15998_),
    .B(_15999_),
    .C(_16001_),
    .Y(_16003_));
 sky130_fd_sc_hd__nand2_1 _38368_ (.A(_16002_),
    .B(_16003_),
    .Y(_16004_));
 sky130_fd_sc_hd__nor2_4 _38369_ (.A(_15785_),
    .B(_15778_),
    .Y(_16005_));
 sky130_fd_sc_hd__nor2_8 _38370_ (.A(_15779_),
    .B(_16005_),
    .Y(_16006_));
 sky130_fd_sc_hd__nand2_1 _38371_ (.A(_16004_),
    .B(_16006_),
    .Y(_16007_));
 sky130_vsdinv _38372_ (.A(_16006_),
    .Y(_16008_));
 sky130_fd_sc_hd__nand3_1 _38373_ (.A(_16002_),
    .B(_16003_),
    .C(_16008_),
    .Y(_16009_));
 sky130_fd_sc_hd__nand2_2 _38374_ (.A(_16007_),
    .B(_16009_),
    .Y(_16010_));
 sky130_fd_sc_hd__nand2_1 _38375_ (.A(_15981_),
    .B(_16010_),
    .Y(_16011_));
 sky130_fd_sc_hd__a21oi_4 _38376_ (.A1(_15998_),
    .A2(_15999_),
    .B1(_16001_),
    .Y(_16012_));
 sky130_fd_sc_hd__nor2_2 _38377_ (.A(_16006_),
    .B(_16012_),
    .Y(_16013_));
 sky130_fd_sc_hd__a21oi_2 _38378_ (.A1(_16002_),
    .A2(_16003_),
    .B1(_16008_),
    .Y(_16014_));
 sky130_fd_sc_hd__a21oi_4 _38379_ (.A1(_16003_),
    .A2(_16013_),
    .B1(_16014_),
    .Y(_16015_));
 sky130_fd_sc_hd__nand3_2 _38380_ (.A(_16015_),
    .B(_15980_),
    .C(_15977_),
    .Y(_16016_));
 sky130_fd_sc_hd__a21oi_4 _38381_ (.A1(_15864_),
    .A2(_15865_),
    .B1(_15862_),
    .Y(_16017_));
 sky130_vsdinv _38382_ (.A(_16017_),
    .Y(_16018_));
 sky130_fd_sc_hd__nand3_4 _38383_ (.A(_16011_),
    .B(_16016_),
    .C(_16018_),
    .Y(_16019_));
 sky130_fd_sc_hd__nand2_1 _38384_ (.A(_15981_),
    .B(_16015_),
    .Y(_16020_));
 sky130_fd_sc_hd__nand3_2 _38385_ (.A(_16010_),
    .B(_15980_),
    .C(_15977_),
    .Y(_16021_));
 sky130_fd_sc_hd__nand3_4 _38386_ (.A(_16020_),
    .B(_16017_),
    .C(_16021_),
    .Y(_16022_));
 sky130_fd_sc_hd__a21boi_4 _38387_ (.A1(_15793_),
    .A2(_15794_),
    .B1_N(_15790_),
    .Y(_16023_));
 sky130_fd_sc_hd__nand2_4 _38388_ (.A(_10990_),
    .B(_11597_),
    .Y(_16024_));
 sky130_fd_sc_hd__nand2_8 _38389_ (.A(_12614_),
    .B(_08616_),
    .Y(_16025_));
 sky130_fd_sc_hd__nor2_8 _38390_ (.A(_16024_),
    .B(_16025_),
    .Y(_16026_));
 sky130_fd_sc_hd__and2_1 _38391_ (.A(_16024_),
    .B(_16025_),
    .X(_16027_));
 sky130_fd_sc_hd__nor2_2 _38392_ (.A(_16026_),
    .B(_16027_),
    .Y(_16028_));
 sky130_fd_sc_hd__or2_4 _38393_ (.A(_15729_),
    .B(_16028_),
    .X(_16029_));
 sky130_fd_sc_hd__nand2_4 _38394_ (.A(_16028_),
    .B(_15729_),
    .Y(_16030_));
 sky130_fd_sc_hd__a2bb2o_2 _38395_ (.A1_N(_15570_),
    .A2_N(_15782_),
    .B1(_15783_),
    .B2(_15781_),
    .X(_16031_));
 sky130_fd_sc_hd__a21oi_4 _38396_ (.A1(_16029_),
    .A2(_16030_),
    .B1(_16031_),
    .Y(_16032_));
 sky130_fd_sc_hd__and3_1 _38397_ (.A(_16029_),
    .B(_16031_),
    .C(_16030_),
    .X(_16033_));
 sky130_fd_sc_hd__nand2_2 _38398_ (.A(_15734_),
    .B(_15732_),
    .Y(_16034_));
 sky130_vsdinv _38399_ (.A(_16034_),
    .Y(_16035_));
 sky130_fd_sc_hd__o21ai_4 _38400_ (.A1(_16032_),
    .A2(_16033_),
    .B1(_16035_),
    .Y(_16036_));
 sky130_fd_sc_hd__nand3_4 _38401_ (.A(_16029_),
    .B(_16031_),
    .C(_16030_),
    .Y(_16037_));
 sky130_fd_sc_hd__nand3b_4 _38402_ (.A_N(_16032_),
    .B(_16034_),
    .C(_16037_),
    .Y(_16038_));
 sky130_fd_sc_hd__nand2_2 _38403_ (.A(_15741_),
    .B(_15738_),
    .Y(_16039_));
 sky130_fd_sc_hd__a21oi_4 _38404_ (.A1(_16036_),
    .A2(_16038_),
    .B1(_16039_),
    .Y(_16040_));
 sky130_fd_sc_hd__nor2_2 _38405_ (.A(_15755_),
    .B(_16040_),
    .Y(_16041_));
 sky130_fd_sc_hd__nand3_2 _38406_ (.A(_16036_),
    .B(_16038_),
    .C(_16039_),
    .Y(_16042_));
 sky130_fd_sc_hd__nand2_1 _38407_ (.A(_16041_),
    .B(_16042_),
    .Y(_16043_));
 sky130_fd_sc_hd__and3_2 _38408_ (.A(_16036_),
    .B(_16038_),
    .C(_16039_),
    .X(_16044_));
 sky130_fd_sc_hd__clkbuf_4 _38409_ (.A(_15754_),
    .X(_16045_));
 sky130_fd_sc_hd__o21ai_2 _38410_ (.A1(_16040_),
    .A2(_16044_),
    .B1(_16045_),
    .Y(_16046_));
 sky130_fd_sc_hd__nand3b_4 _38411_ (.A_N(_16023_),
    .B(_16043_),
    .C(_16046_),
    .Y(_16047_));
 sky130_fd_sc_hd__buf_4 _38412_ (.A(_15748_),
    .X(_16048_));
 sky130_fd_sc_hd__o21ai_2 _38413_ (.A1(_16040_),
    .A2(_16044_),
    .B1(_16048_),
    .Y(_16049_));
 sky130_fd_sc_hd__nand3b_2 _38414_ (.A_N(_16040_),
    .B(_16045_),
    .C(_16042_),
    .Y(_16050_));
 sky130_fd_sc_hd__nand3_4 _38415_ (.A(_16049_),
    .B(_16050_),
    .C(_16023_),
    .Y(_16051_));
 sky130_fd_sc_hd__nor2_1 _38416_ (.A(_15755_),
    .B(_15750_),
    .Y(_16052_));
 sky130_fd_sc_hd__nor2_2 _38417_ (.A(_15752_),
    .B(_16052_),
    .Y(_16053_));
 sky130_vsdinv _38418_ (.A(_16053_),
    .Y(_16054_));
 sky130_fd_sc_hd__a21oi_4 _38419_ (.A1(_16047_),
    .A2(_16051_),
    .B1(_16054_),
    .Y(_16055_));
 sky130_fd_sc_hd__nand2_1 _38420_ (.A(_16047_),
    .B(_16051_),
    .Y(_16056_));
 sky130_fd_sc_hd__nor2_1 _38421_ (.A(_16053_),
    .B(_16056_),
    .Y(_16057_));
 sky130_fd_sc_hd__o2bb2ai_2 _38422_ (.A1_N(_16019_),
    .A2_N(_16022_),
    .B1(_16055_),
    .B2(_16057_),
    .Y(_16058_));
 sky130_fd_sc_hd__and2_1 _38423_ (.A(_16051_),
    .B(_16054_),
    .X(_16059_));
 sky130_fd_sc_hd__a21oi_4 _38424_ (.A1(_16059_),
    .A2(_16047_),
    .B1(_16055_),
    .Y(_16060_));
 sky130_fd_sc_hd__nand3_4 _38425_ (.A(_16060_),
    .B(_16019_),
    .C(_16022_),
    .Y(_16061_));
 sky130_fd_sc_hd__nand2_1 _38426_ (.A(_16058_),
    .B(_16061_),
    .Y(_16062_));
 sky130_fd_sc_hd__nand2_2 _38427_ (.A(_15880_),
    .B(_15879_),
    .Y(_16063_));
 sky130_vsdinv _38428_ (.A(_16063_),
    .Y(_16064_));
 sky130_fd_sc_hd__nand2_4 _38429_ (.A(_16062_),
    .B(_16064_),
    .Y(_16065_));
 sky130_fd_sc_hd__nand3_4 _38430_ (.A(_16058_),
    .B(_16061_),
    .C(_16063_),
    .Y(_16066_));
 sky130_fd_sc_hd__nor2_8 _38431_ (.A(_15697_),
    .B(_15746_),
    .Y(_16067_));
 sky130_fd_sc_hd__a31o_1 _38432_ (.A1(_15471_),
    .A2(_15705_),
    .A3(_15703_),
    .B1(_15699_),
    .X(_16068_));
 sky130_fd_sc_hd__nor2_1 _38433_ (.A(_16067_),
    .B(_16068_),
    .Y(_16069_));
 sky130_fd_sc_hd__nand2_1 _38434_ (.A(_16068_),
    .B(_16067_),
    .Y(_16070_));
 sky130_fd_sc_hd__or2b_1 _38435_ (.A(_16069_),
    .B_N(_16070_),
    .X(_16071_));
 sky130_fd_sc_hd__nand2_1 _38436_ (.A(_16071_),
    .B(_14283_),
    .Y(_16072_));
 sky130_vsdinv _38437_ (.A(_16069_),
    .Y(_16073_));
 sky130_fd_sc_hd__nand3_1 _38438_ (.A(_16073_),
    .B(_13989_),
    .C(_16070_),
    .Y(_16074_));
 sky130_fd_sc_hd__nand2_1 _38439_ (.A(_16072_),
    .B(_16074_),
    .Y(_16075_));
 sky130_fd_sc_hd__or2b_1 _38440_ (.A(_15877_),
    .B_N(_15757_),
    .X(_16076_));
 sky130_fd_sc_hd__nor2_1 _38441_ (.A(_16075_),
    .B(_16076_),
    .Y(_16077_));
 sky130_fd_sc_hd__nand2_2 _38442_ (.A(_16076_),
    .B(_16075_),
    .Y(_16078_));
 sky130_fd_sc_hd__or2b_1 _38443_ (.A(_16077_),
    .B_N(_16078_),
    .X(_16079_));
 sky130_fd_sc_hd__nand2_2 _38444_ (.A(_15712_),
    .B(_15710_),
    .Y(_16080_));
 sky130_fd_sc_hd__nand2_1 _38445_ (.A(_16079_),
    .B(_16080_),
    .Y(_16081_));
 sky130_fd_sc_hd__and2b_1 _38446_ (.A_N(_16077_),
    .B(_16078_),
    .X(_16082_));
 sky130_vsdinv _38447_ (.A(_16080_),
    .Y(_16083_));
 sky130_fd_sc_hd__nand2_1 _38448_ (.A(_16082_),
    .B(_16083_),
    .Y(_16084_));
 sky130_fd_sc_hd__nand2_2 _38449_ (.A(_16081_),
    .B(_16084_),
    .Y(_16085_));
 sky130_fd_sc_hd__a21o_1 _38450_ (.A1(_16065_),
    .A2(_16066_),
    .B1(_16085_),
    .X(_16086_));
 sky130_fd_sc_hd__nand2_1 _38451_ (.A(_15888_),
    .B(_15891_),
    .Y(_16087_));
 sky130_fd_sc_hd__nand2_2 _38452_ (.A(_16087_),
    .B(_15892_),
    .Y(_16088_));
 sky130_fd_sc_hd__nand3_2 _38453_ (.A(_16065_),
    .B(_16085_),
    .C(_16066_),
    .Y(_16089_));
 sky130_fd_sc_hd__nand3_4 _38454_ (.A(_16086_),
    .B(_16088_),
    .C(_16089_),
    .Y(_16090_));
 sky130_fd_sc_hd__nor2_1 _38455_ (.A(_16083_),
    .B(_16082_),
    .Y(_16091_));
 sky130_vsdinv _38456_ (.A(_16084_),
    .Y(_16092_));
 sky130_fd_sc_hd__o2bb2ai_2 _38457_ (.A1_N(_16066_),
    .A2_N(_16065_),
    .B1(_16091_),
    .B2(_16092_),
    .Y(_16093_));
 sky130_fd_sc_hd__nand2_1 _38458_ (.A(_16079_),
    .B(_16083_),
    .Y(_16094_));
 sky130_fd_sc_hd__nand2_2 _38459_ (.A(_16082_),
    .B(_16080_),
    .Y(_16095_));
 sky130_fd_sc_hd__nand2_2 _38460_ (.A(_16094_),
    .B(_16095_),
    .Y(_16096_));
 sky130_fd_sc_hd__nand3_4 _38461_ (.A(_16065_),
    .B(_16096_),
    .C(_16066_),
    .Y(_16097_));
 sky130_fd_sc_hd__nand3b_4 _38462_ (.A_N(_16088_),
    .B(_16093_),
    .C(_16097_),
    .Y(_16098_));
 sky130_fd_sc_hd__and3_2 _38463_ (.A(_15721_),
    .B(_14329_),
    .C(_15720_),
    .X(_16099_));
 sky130_fd_sc_hd__nor2_2 _38464_ (.A(_15889_),
    .B(_15722_),
    .Y(_16100_));
 sky130_fd_sc_hd__nor2_4 _38465_ (.A(_14330_),
    .B(_16100_),
    .Y(_16101_));
 sky130_fd_sc_hd__nor2_4 _38466_ (.A(_16099_),
    .B(_16101_),
    .Y(_16102_));
 sky130_vsdinv _38467_ (.A(_16102_),
    .Y(_16103_));
 sky130_fd_sc_hd__a21o_1 _38468_ (.A1(_16090_),
    .A2(_16098_),
    .B1(_16103_),
    .X(_16104_));
 sky130_fd_sc_hd__a21boi_4 _38469_ (.A1(_15898_),
    .A2(_15906_),
    .B1_N(_15894_),
    .Y(_16105_));
 sky130_fd_sc_hd__nand3_4 _38470_ (.A(_16090_),
    .B(_16098_),
    .C(_16103_),
    .Y(_16106_));
 sky130_fd_sc_hd__nand3_2 _38471_ (.A(_16104_),
    .B(_16105_),
    .C(_16106_),
    .Y(_16107_));
 sky130_fd_sc_hd__o2bb2ai_2 _38472_ (.A1_N(_16098_),
    .A2_N(_16090_),
    .B1(_16101_),
    .B2(_16099_),
    .Y(_16108_));
 sky130_fd_sc_hd__nand3_4 _38473_ (.A(_16090_),
    .B(_16098_),
    .C(_16102_),
    .Y(_16109_));
 sky130_fd_sc_hd__nand3b_4 _38474_ (.A_N(_16105_),
    .B(_16108_),
    .C(_16109_),
    .Y(_16110_));
 sky130_fd_sc_hd__a21oi_1 _38475_ (.A1(_16107_),
    .A2(_16110_),
    .B1(_15901_),
    .Y(_16111_));
 sky130_fd_sc_hd__a21oi_4 _38476_ (.A1(_16104_),
    .A2(_16106_),
    .B1(_16105_),
    .Y(_16112_));
 sky130_fd_sc_hd__nand2_2 _38477_ (.A(_16107_),
    .B(_15901_),
    .Y(_16113_));
 sky130_fd_sc_hd__nor2_1 _38478_ (.A(_16112_),
    .B(_16113_),
    .Y(_16114_));
 sky130_fd_sc_hd__a21bo_1 _38479_ (.A1(_15665_),
    .A2(_15914_),
    .B1_N(_15908_),
    .X(_16115_));
 sky130_fd_sc_hd__o21bai_2 _38480_ (.A1(_16111_),
    .A2(_16114_),
    .B1_N(_16115_),
    .Y(_16116_));
 sky130_fd_sc_hd__a21o_1 _38481_ (.A1(_16107_),
    .A2(_16110_),
    .B1(_15901_),
    .X(_16117_));
 sky130_fd_sc_hd__o211ai_4 _38482_ (.A1(_16112_),
    .A2(_16113_),
    .B1(_16115_),
    .C1(_16117_),
    .Y(_16118_));
 sky130_fd_sc_hd__and2_1 _38483_ (.A(_16116_),
    .B(_16118_),
    .X(_16119_));
 sky130_vsdinv _38484_ (.A(_15435_),
    .Y(_16120_));
 sky130_fd_sc_hd__o2bb2ai_2 _38485_ (.A1_N(_15431_),
    .A2_N(_15429_),
    .B1(_15191_),
    .B2(_15434_),
    .Y(_16121_));
 sky130_fd_sc_hd__o2111ai_4 _38486_ (.A1(_16120_),
    .A2(_16121_),
    .B1(_15183_),
    .C1(_15433_),
    .D1(_15178_),
    .Y(_16122_));
 sky130_fd_sc_hd__o2111ai_4 _38487_ (.A1(_15679_),
    .A2(_15685_),
    .B1(_15922_),
    .C1(_15687_),
    .D1(_15919_),
    .Y(_16123_));
 sky130_fd_sc_hd__nor2_8 _38488_ (.A(_16122_),
    .B(_16123_),
    .Y(_16124_));
 sky130_fd_sc_hd__and4_1 _38489_ (.A(_14338_),
    .B(_14023_),
    .C(_14024_),
    .D(_14339_),
    .X(_16125_));
 sky130_fd_sc_hd__nand3_2 _38490_ (.A(_16124_),
    .B(_16125_),
    .C(_15185_),
    .Y(_16126_));
 sky130_fd_sc_hd__a21boi_2 _38491_ (.A1(_15694_),
    .A2(_15919_),
    .B1_N(_15922_),
    .Y(_16127_));
 sky130_fd_sc_hd__o21ai_4 _38492_ (.A1(_15692_),
    .A2(_16123_),
    .B1(_16127_),
    .Y(_16128_));
 sky130_fd_sc_hd__a21oi_1 _38493_ (.A1(_15189_),
    .A2(_16124_),
    .B1(_16128_),
    .Y(_16129_));
 sky130_fd_sc_hd__o21a_4 _38494_ (.A1(_16126_),
    .A2(_14032_),
    .B1(_16129_),
    .X(_16130_));
 sky130_fd_sc_hd__nand3_4 _38495_ (.A(_15690_),
    .B(_15688_),
    .C(_15923_),
    .Y(_16131_));
 sky130_fd_sc_hd__nand3_1 _38496_ (.A(_14340_),
    .B(_14025_),
    .C(_15185_),
    .Y(_16132_));
 sky130_fd_sc_hd__nor2_2 _38497_ (.A(_16131_),
    .B(_16132_),
    .Y(_16133_));
 sky130_fd_sc_hd__nand3_4 _38498_ (.A(net409),
    .B(_14029_),
    .C(_16133_),
    .Y(_16134_));
 sky130_fd_sc_hd__nand2_2 _38499_ (.A(_16130_),
    .B(_16134_),
    .Y(_16135_));
 sky130_fd_sc_hd__or2_1 _38500_ (.A(_16119_),
    .B(_16135_),
    .X(_16136_));
 sky130_fd_sc_hd__nand2_1 _38501_ (.A(_16135_),
    .B(_16119_),
    .Y(_16137_));
 sky130_fd_sc_hd__and2_2 _38502_ (.A(_16136_),
    .B(_16137_),
    .X(_02667_));
 sky130_fd_sc_hd__a21boi_2 _38503_ (.A1(_16093_),
    .A2(_16097_),
    .B1_N(_16088_),
    .Y(_16138_));
 sky130_fd_sc_hd__a21o_1 _38504_ (.A1(_16098_),
    .A2(_16102_),
    .B1(_16138_),
    .X(_16139_));
 sky130_fd_sc_hd__nand2_2 _38505_ (.A(_16051_),
    .B(_16054_),
    .Y(_16140_));
 sky130_fd_sc_hd__nor2_8 _38506_ (.A(_15704_),
    .B(_16067_),
    .Y(_16141_));
 sky130_vsdinv _38507_ (.A(_16141_),
    .Y(_16142_));
 sky130_fd_sc_hd__nand2_2 _38508_ (.A(_16067_),
    .B(_15700_),
    .Y(_16143_));
 sky130_fd_sc_hd__and3_1 _38509_ (.A(_13654_),
    .B(_16142_),
    .C(_16143_),
    .X(_16144_));
 sky130_vsdinv _38510_ (.A(_16143_),
    .Y(_16145_));
 sky130_fd_sc_hd__o21ai_1 _38511_ (.A1(_16141_),
    .A2(_16145_),
    .B1(_13655_),
    .Y(_16146_));
 sky130_fd_sc_hd__and2b_1 _38512_ (.A_N(_16144_),
    .B(_16146_),
    .X(_16147_));
 sky130_vsdinv _38513_ (.A(_16147_),
    .Y(_16148_));
 sky130_fd_sc_hd__buf_4 _38514_ (.A(_16148_),
    .X(_16149_));
 sky130_fd_sc_hd__a21o_1 _38515_ (.A1(_16140_),
    .A2(_16047_),
    .B1(_16149_),
    .X(_16150_));
 sky130_fd_sc_hd__nand3_4 _38516_ (.A(_16149_),
    .B(_16047_),
    .C(_16140_),
    .Y(_16151_));
 sky130_fd_sc_hd__nand2_1 _38517_ (.A(_16150_),
    .B(_16151_),
    .Y(_16152_));
 sky130_fd_sc_hd__a21oi_2 _38518_ (.A1(_16071_),
    .A2(_13989_),
    .B1(_16141_),
    .Y(_16153_));
 sky130_fd_sc_hd__and2_1 _38519_ (.A(_16152_),
    .B(_16153_),
    .X(_16154_));
 sky130_fd_sc_hd__nand3b_4 _38520_ (.A_N(_16153_),
    .B(_16150_),
    .C(_16151_),
    .Y(_16155_));
 sky130_vsdinv _38521_ (.A(_16155_),
    .Y(_16156_));
 sky130_fd_sc_hd__nand2_2 _38522_ (.A(_15950_),
    .B(_15946_),
    .Y(_16157_));
 sky130_fd_sc_hd__nand2_2 _38523_ (.A(_19593_),
    .B(_19864_),
    .Y(_16158_));
 sky130_fd_sc_hd__buf_2 _38524_ (.A(_15931_),
    .X(_16159_));
 sky130_fd_sc_hd__o22a_2 _38525_ (.A1(_16159_),
    .A2(_08080_),
    .B1(_15932_),
    .B2(_12916_),
    .X(_16160_));
 sky130_fd_sc_hd__a311o_1 _38526_ (.A1(_19867_),
    .A2(_15930_),
    .A3(_19870_),
    .B1(_16158_),
    .C1(_16160_),
    .X(_16161_));
 sky130_fd_sc_hd__and3_1 _38527_ (.A(_15929_),
    .B(_19867_),
    .C(_11724_),
    .X(_16162_));
 sky130_fd_sc_hd__o21ai_1 _38528_ (.A1(_16160_),
    .A2(_16162_),
    .B1(_16158_),
    .Y(_16163_));
 sky130_fd_sc_hd__nand2_1 _38529_ (.A(_16161_),
    .B(_16163_),
    .Y(_16164_));
 sky130_vsdinv _38530_ (.A(_16164_),
    .Y(_16165_));
 sky130_fd_sc_hd__and4_2 _38531_ (.A(_08447_),
    .B(_15937_),
    .C(_19577_),
    .D(_14452_),
    .X(_16166_));
 sky130_fd_sc_hd__o22a_2 _38532_ (.A1(_19879_),
    .A2(_18475_),
    .B1(_15939_),
    .B2(_10732_),
    .X(_16167_));
 sky130_fd_sc_hd__nor2_1 _38533_ (.A(_16166_),
    .B(_16167_),
    .Y(_16168_));
 sky130_fd_sc_hd__nor2_2 _38534_ (.A(_15823_),
    .B(_10971_),
    .Y(_16169_));
 sky130_fd_sc_hd__nand2_2 _38535_ (.A(_16168_),
    .B(_16169_),
    .Y(_16170_));
 sky130_fd_sc_hd__o21bai_2 _38536_ (.A1(_16166_),
    .A2(_16167_),
    .B1_N(_16169_),
    .Y(_16171_));
 sky130_fd_sc_hd__nand2_1 _38537_ (.A(_16170_),
    .B(_16171_),
    .Y(_16172_));
 sky130_fd_sc_hd__nor2_2 _38538_ (.A(_15943_),
    .B(_15940_),
    .Y(_16173_));
 sky130_fd_sc_hd__nor2_4 _38539_ (.A(_15938_),
    .B(_16173_),
    .Y(_16174_));
 sky130_fd_sc_hd__nand2_2 _38540_ (.A(_16172_),
    .B(_16174_),
    .Y(_16175_));
 sky130_fd_sc_hd__nand3b_4 _38541_ (.A_N(_16174_),
    .B(_16170_),
    .C(_16171_),
    .Y(_16176_));
 sky130_fd_sc_hd__nand3_4 _38542_ (.A(_16165_),
    .B(_16175_),
    .C(_16176_),
    .Y(_16177_));
 sky130_fd_sc_hd__nand2_1 _38543_ (.A(_16176_),
    .B(_16175_),
    .Y(_16178_));
 sky130_fd_sc_hd__nand2_2 _38544_ (.A(_16178_),
    .B(_16164_),
    .Y(_16179_));
 sky130_fd_sc_hd__nand3_4 _38545_ (.A(_16157_),
    .B(_16177_),
    .C(_16179_),
    .Y(_16180_));
 sky130_fd_sc_hd__nand2_1 _38546_ (.A(_16179_),
    .B(_16177_),
    .Y(_16181_));
 sky130_fd_sc_hd__nand3_4 _38547_ (.A(_16181_),
    .B(_15946_),
    .C(_15950_),
    .Y(_16182_));
 sky130_fd_sc_hd__and4_4 _38548_ (.A(_19598_),
    .B(_19601_),
    .C(_14501_),
    .D(_13413_),
    .X(_16183_));
 sky130_fd_sc_hd__buf_2 _38549_ (.A(_15957_),
    .X(_16184_));
 sky130_fd_sc_hd__o22a_2 _38550_ (.A1(_15956_),
    .A2(_15802_),
    .B1(_16184_),
    .B2(_10652_),
    .X(_16185_));
 sky130_fd_sc_hd__nor2_1 _38551_ (.A(_08579_),
    .B(_13855_),
    .Y(_16186_));
 sky130_vsdinv _38552_ (.A(_16186_),
    .Y(_16187_));
 sky130_fd_sc_hd__nor3_4 _38553_ (.A(_16183_),
    .B(_16185_),
    .C(_16187_),
    .Y(_16188_));
 sky130_vsdinv _38554_ (.A(_16188_),
    .Y(_16189_));
 sky130_fd_sc_hd__o21ai_2 _38555_ (.A1(_16183_),
    .A2(_16185_),
    .B1(_16187_),
    .Y(_16190_));
 sky130_fd_sc_hd__o32a_2 _38556_ (.A1(_08080_),
    .A2(_10971_),
    .A3(_15928_),
    .B1(_15927_),
    .B2(_15933_),
    .X(_16191_));
 sky130_fd_sc_hd__a21boi_2 _38557_ (.A1(_16189_),
    .A2(_16190_),
    .B1_N(_16191_),
    .Y(_16192_));
 sky130_fd_sc_hd__nand2_1 _38558_ (.A(_16189_),
    .B(_16190_),
    .Y(_16193_));
 sky130_fd_sc_hd__nor2_1 _38559_ (.A(_16191_),
    .B(_16193_),
    .Y(_16194_));
 sky130_vsdinv _38560_ (.A(_15955_),
    .Y(_16195_));
 sky130_fd_sc_hd__and2_1 _38561_ (.A(_15959_),
    .B(_16195_),
    .X(_16196_));
 sky130_fd_sc_hd__o21ai_2 _38562_ (.A1(_16192_),
    .A2(_16194_),
    .B1(_16196_),
    .Y(_16197_));
 sky130_vsdinv _38563_ (.A(_16197_),
    .Y(_16198_));
 sky130_fd_sc_hd__or3b_4 _38564_ (.A(_16188_),
    .B(_16191_),
    .C_N(_16190_),
    .X(_16199_));
 sky130_fd_sc_hd__nand2_1 _38565_ (.A(_15959_),
    .B(_16195_),
    .Y(_16200_));
 sky130_fd_sc_hd__nand2_1 _38566_ (.A(_16193_),
    .B(_16191_),
    .Y(_16201_));
 sky130_fd_sc_hd__nand3_2 _38567_ (.A(_16199_),
    .B(_16200_),
    .C(_16201_),
    .Y(_16202_));
 sky130_vsdinv _38568_ (.A(_16202_),
    .Y(_16203_));
 sky130_fd_sc_hd__o2bb2ai_4 _38569_ (.A1_N(_16180_),
    .A2_N(_16182_),
    .B1(_16198_),
    .B2(_16203_),
    .Y(_16204_));
 sky130_fd_sc_hd__nand2_2 _38570_ (.A(_16197_),
    .B(_16202_),
    .Y(_16205_));
 sky130_fd_sc_hd__nand3b_4 _38571_ (.A_N(_16205_),
    .B(_16180_),
    .C(_16182_),
    .Y(_16206_));
 sky130_fd_sc_hd__o21ai_4 _38572_ (.A1(_15952_),
    .A2(_15975_),
    .B1(_15973_),
    .Y(_16207_));
 sky130_fd_sc_hd__a21oi_4 _38573_ (.A1(_16204_),
    .A2(_16206_),
    .B1(_16207_),
    .Y(_16208_));
 sky130_vsdinv _38574_ (.A(_16180_),
    .Y(_16209_));
 sky130_fd_sc_hd__nand3_1 _38575_ (.A(_16182_),
    .B(_16197_),
    .C(_16202_),
    .Y(_16210_));
 sky130_fd_sc_hd__o211a_2 _38576_ (.A1(_16209_),
    .A2(_16210_),
    .B1(_16204_),
    .C1(_16207_),
    .X(_16211_));
 sky130_fd_sc_hd__nor2_2 _38577_ (.A(_15962_),
    .B(_15961_),
    .Y(_16212_));
 sky130_fd_sc_hd__a21o_1 _38578_ (.A1(_15963_),
    .A2(_15965_),
    .B1(_16212_),
    .X(_16213_));
 sky130_fd_sc_hd__nand2_2 _38579_ (.A(_19608_),
    .B(_11909_),
    .Y(_16214_));
 sky130_fd_sc_hd__nand2_2 _38580_ (.A(_12466_),
    .B(_11178_),
    .Y(_16215_));
 sky130_fd_sc_hd__or2_2 _38581_ (.A(_16214_),
    .B(_16215_),
    .X(_16216_));
 sky130_fd_sc_hd__nand2_2 _38582_ (.A(_16214_),
    .B(_16215_),
    .Y(_16217_));
 sky130_fd_sc_hd__nand2_1 _38583_ (.A(_19618_),
    .B(_11583_),
    .Y(_16218_));
 sky130_fd_sc_hd__a21bo_1 _38584_ (.A1(_16216_),
    .A2(_16217_),
    .B1_N(_16218_),
    .X(_16219_));
 sky130_fd_sc_hd__nand3b_4 _38585_ (.A_N(_16218_),
    .B(_16216_),
    .C(_16217_),
    .Y(_16220_));
 sky130_fd_sc_hd__a31o_1 _38586_ (.A1(_15984_),
    .A2(_19619_),
    .A3(_19846_),
    .B1(_15982_),
    .X(_16221_));
 sky130_fd_sc_hd__a21o_1 _38587_ (.A1(_16219_),
    .A2(_16220_),
    .B1(_16221_),
    .X(_16222_));
 sky130_fd_sc_hd__nand3_4 _38588_ (.A(_16219_),
    .B(_16221_),
    .C(_16220_),
    .Y(_16223_));
 sky130_fd_sc_hd__nand2_1 _38589_ (.A(_19629_),
    .B(_19827_),
    .Y(_16224_));
 sky130_fd_sc_hd__nand2_4 _38590_ (.A(_19622_),
    .B(_11202_),
    .Y(_16225_));
 sky130_fd_sc_hd__nand2_2 _38591_ (.A(_19623_),
    .B(_19835_),
    .Y(_16226_));
 sky130_fd_sc_hd__o21ai_1 _38592_ (.A1(_15993_),
    .A2(_10597_),
    .B1(_16226_),
    .Y(_16227_));
 sky130_fd_sc_hd__o21ai_2 _38593_ (.A1(_15995_),
    .A2(_16225_),
    .B1(_16227_),
    .Y(_16228_));
 sky130_fd_sc_hd__nor2_4 _38594_ (.A(_16224_),
    .B(_16228_),
    .Y(_16229_));
 sky130_fd_sc_hd__and2_1 _38595_ (.A(_16228_),
    .B(_16224_),
    .X(_16230_));
 sky130_fd_sc_hd__nor2_2 _38596_ (.A(_16229_),
    .B(_16230_),
    .Y(_16231_));
 sky130_fd_sc_hd__a21o_1 _38597_ (.A1(_16222_),
    .A2(_16223_),
    .B1(_16231_),
    .X(_16232_));
 sky130_fd_sc_hd__nand3_4 _38598_ (.A(_16222_),
    .B(_16223_),
    .C(_16231_),
    .Y(_16233_));
 sky130_fd_sc_hd__nand3_4 _38599_ (.A(_16213_),
    .B(_16232_),
    .C(_16233_),
    .Y(_16234_));
 sky130_fd_sc_hd__nand2_2 _38600_ (.A(_16232_),
    .B(_16233_),
    .Y(_16235_));
 sky130_fd_sc_hd__a21oi_4 _38601_ (.A1(_15963_),
    .A2(_15965_),
    .B1(_16212_),
    .Y(_16236_));
 sky130_fd_sc_hd__nand2_2 _38602_ (.A(_16235_),
    .B(_16236_),
    .Y(_16237_));
 sky130_fd_sc_hd__nand2_2 _38603_ (.A(_15999_),
    .B(_15990_),
    .Y(_16238_));
 sky130_fd_sc_hd__a21o_1 _38604_ (.A1(_16234_),
    .A2(_16237_),
    .B1(_16238_),
    .X(_16239_));
 sky130_fd_sc_hd__nand3_4 _38605_ (.A(_16234_),
    .B(_16238_),
    .C(_16237_),
    .Y(_16240_));
 sky130_fd_sc_hd__and2_2 _38606_ (.A(_16239_),
    .B(_16240_),
    .X(_16241_));
 sky130_fd_sc_hd__o21ai_2 _38607_ (.A1(_16208_),
    .A2(_16211_),
    .B1(_16241_),
    .Y(_16242_));
 sky130_fd_sc_hd__a21boi_4 _38608_ (.A1(_16015_),
    .A2(_15977_),
    .B1_N(_15980_),
    .Y(_16243_));
 sky130_fd_sc_hd__a21o_2 _38609_ (.A1(_16204_),
    .A2(_16206_),
    .B1(_16207_),
    .X(_16244_));
 sky130_fd_sc_hd__nand3_4 _38610_ (.A(_16207_),
    .B(_16204_),
    .C(_16206_),
    .Y(_16245_));
 sky130_fd_sc_hd__nand2_4 _38611_ (.A(_16239_),
    .B(_16240_),
    .Y(_16246_));
 sky130_fd_sc_hd__nand3_4 _38612_ (.A(_16244_),
    .B(_16245_),
    .C(_16246_),
    .Y(_16247_));
 sky130_fd_sc_hd__nand3_4 _38613_ (.A(_16242_),
    .B(_16243_),
    .C(_16247_),
    .Y(_16248_));
 sky130_fd_sc_hd__o21ai_2 _38614_ (.A1(_16208_),
    .A2(_16211_),
    .B1(_16246_),
    .Y(_16249_));
 sky130_fd_sc_hd__a21oi_2 _38615_ (.A1(_15978_),
    .A2(_15979_),
    .B1(_15970_),
    .Y(_16250_));
 sky130_fd_sc_hd__o21ai_2 _38616_ (.A1(_16010_),
    .A2(_16250_),
    .B1(_15980_),
    .Y(_16251_));
 sky130_fd_sc_hd__nand3_4 _38617_ (.A(_16244_),
    .B(_16241_),
    .C(_16245_),
    .Y(_16252_));
 sky130_fd_sc_hd__nand3_4 _38618_ (.A(_16249_),
    .B(_16251_),
    .C(_16252_),
    .Y(_16253_));
 sky130_fd_sc_hd__o21ai_2 _38619_ (.A1(_16035_),
    .A2(_16032_),
    .B1(_16037_),
    .Y(_16254_));
 sky130_fd_sc_hd__o32a_1 _38620_ (.A1(_15993_),
    .A2(_12902_),
    .A3(_16226_),
    .B1(_15991_),
    .B2(_15996_),
    .X(_16255_));
 sky130_vsdinv _38621_ (.A(_10998_),
    .Y(_16256_));
 sky130_fd_sc_hd__nor2_4 _38622_ (.A(_16025_),
    .B(_16256_),
    .Y(_16257_));
 sky130_fd_sc_hd__o21a_4 _38623_ (.A1(_08615_),
    .A2(_08616_),
    .B1(_11593_),
    .X(_16258_));
 sky130_fd_sc_hd__nand2_2 _38624_ (.A(_16258_),
    .B(_19642_),
    .Y(_16259_));
 sky130_fd_sc_hd__or2_2 _38625_ (.A(_16257_),
    .B(_16259_),
    .X(_16260_));
 sky130_vsdinv _38626_ (.A(_16258_),
    .Y(_16261_));
 sky130_fd_sc_hd__o21ai_2 _38627_ (.A1(_16257_),
    .A2(_16261_),
    .B1(_15730_),
    .Y(_16262_));
 sky130_fd_sc_hd__nand2_2 _38628_ (.A(_16260_),
    .B(_16262_),
    .Y(_16263_));
 sky130_fd_sc_hd__nand2_2 _38629_ (.A(_16255_),
    .B(_16263_),
    .Y(_16264_));
 sky130_fd_sc_hd__and2_4 _38630_ (.A(_16260_),
    .B(_16262_),
    .X(_16265_));
 sky130_fd_sc_hd__o32ai_4 _38631_ (.A1(_15993_),
    .A2(_12902_),
    .A3(_16226_),
    .B1(_15991_),
    .B2(_15996_),
    .Y(_16266_));
 sky130_fd_sc_hd__nand2_4 _38632_ (.A(_16265_),
    .B(_16266_),
    .Y(_16267_));
 sky130_fd_sc_hd__nand2_1 _38633_ (.A(_16264_),
    .B(_16267_),
    .Y(_16268_));
 sky130_vsdinv _38634_ (.A(_16030_),
    .Y(_16269_));
 sky130_fd_sc_hd__nor2_8 _38635_ (.A(_16026_),
    .B(_16269_),
    .Y(_16270_));
 sky130_vsdinv _38636_ (.A(_16270_),
    .Y(_16271_));
 sky130_fd_sc_hd__nand2_1 _38637_ (.A(_16268_),
    .B(_16271_),
    .Y(_16272_));
 sky130_fd_sc_hd__nand3_2 _38638_ (.A(_16264_),
    .B(_16267_),
    .C(_16270_),
    .Y(_16273_));
 sky130_fd_sc_hd__nand3b_4 _38639_ (.A_N(_16254_),
    .B(_16272_),
    .C(_16273_),
    .Y(_16274_));
 sky130_fd_sc_hd__nand2_1 _38640_ (.A(_16268_),
    .B(_16270_),
    .Y(_16275_));
 sky130_fd_sc_hd__nand3_2 _38641_ (.A(_16271_),
    .B(_16264_),
    .C(_16267_),
    .Y(_16276_));
 sky130_fd_sc_hd__nand3_4 _38642_ (.A(_16275_),
    .B(_16254_),
    .C(_16276_),
    .Y(_16277_));
 sky130_fd_sc_hd__nand3_2 _38643_ (.A(_16274_),
    .B(_16277_),
    .C(_15755_),
    .Y(_16278_));
 sky130_fd_sc_hd__nand2_1 _38644_ (.A(_16274_),
    .B(_16277_),
    .Y(_16279_));
 sky130_fd_sc_hd__nand2_1 _38645_ (.A(_16279_),
    .B(_16048_),
    .Y(_16280_));
 sky130_fd_sc_hd__o2111ai_4 _38646_ (.A1(_16012_),
    .A2(_16006_),
    .B1(_16003_),
    .C1(_16278_),
    .D1(_16280_),
    .Y(_16281_));
 sky130_fd_sc_hd__o21ai_2 _38647_ (.A1(_16006_),
    .A2(_16012_),
    .B1(_16003_),
    .Y(_16282_));
 sky130_fd_sc_hd__nand2_1 _38648_ (.A(_16279_),
    .B(_16045_),
    .Y(_16283_));
 sky130_fd_sc_hd__nand3_2 _38649_ (.A(_16274_),
    .B(_16277_),
    .C(_15758_),
    .Y(_16284_));
 sky130_fd_sc_hd__nand3_4 _38650_ (.A(_16282_),
    .B(_16283_),
    .C(_16284_),
    .Y(_16285_));
 sky130_fd_sc_hd__nor2_4 _38651_ (.A(_16044_),
    .B(_16041_),
    .Y(_16286_));
 sky130_fd_sc_hd__a21boi_4 _38652_ (.A1(_16281_),
    .A2(_16285_),
    .B1_N(_16286_),
    .Y(_16287_));
 sky130_fd_sc_hd__nand2_2 _38653_ (.A(_16281_),
    .B(_16285_),
    .Y(_16288_));
 sky130_fd_sc_hd__nor2_4 _38654_ (.A(_16286_),
    .B(_16288_),
    .Y(_16289_));
 sky130_fd_sc_hd__o2bb2ai_4 _38655_ (.A1_N(_16248_),
    .A2_N(_16253_),
    .B1(_16287_),
    .B2(_16289_),
    .Y(_16290_));
 sky130_fd_sc_hd__nor2_2 _38656_ (.A(_16287_),
    .B(_16289_),
    .Y(_16291_));
 sky130_fd_sc_hd__nand3_4 _38657_ (.A(_16291_),
    .B(_16253_),
    .C(_16248_),
    .Y(_16292_));
 sky130_fd_sc_hd__nand2_1 _38658_ (.A(_16060_),
    .B(_16022_),
    .Y(_16293_));
 sky130_fd_sc_hd__nand2_4 _38659_ (.A(_16293_),
    .B(_16019_),
    .Y(_16294_));
 sky130_fd_sc_hd__a21oi_4 _38660_ (.A1(_16290_),
    .A2(_16292_),
    .B1(_16294_),
    .Y(_16295_));
 sky130_fd_sc_hd__and3_1 _38661_ (.A(_16249_),
    .B(_16251_),
    .C(_16252_),
    .X(_16296_));
 sky130_fd_sc_hd__nand2_1 _38662_ (.A(_16291_),
    .B(_16248_),
    .Y(_16297_));
 sky130_fd_sc_hd__o211a_1 _38663_ (.A1(_16296_),
    .A2(_16297_),
    .B1(_16290_),
    .C1(_16294_),
    .X(_16298_));
 sky130_fd_sc_hd__o22ai_4 _38664_ (.A1(_16154_),
    .A2(_16156_),
    .B1(_16295_),
    .B2(_16298_),
    .Y(_16299_));
 sky130_fd_sc_hd__a21oi_1 _38665_ (.A1(_16058_),
    .A2(_16061_),
    .B1(_16063_),
    .Y(_16300_));
 sky130_fd_sc_hd__o21ai_2 _38666_ (.A1(_16300_),
    .A2(_16096_),
    .B1(_16066_),
    .Y(_16301_));
 sky130_fd_sc_hd__a21o_1 _38667_ (.A1(_16290_),
    .A2(_16292_),
    .B1(_16294_),
    .X(_16302_));
 sky130_fd_sc_hd__nand2_1 _38668_ (.A(_16152_),
    .B(_16153_),
    .Y(_16303_));
 sky130_fd_sc_hd__nand2_2 _38669_ (.A(_16303_),
    .B(_16155_),
    .Y(_16304_));
 sky130_vsdinv _38670_ (.A(_16304_),
    .Y(_16305_));
 sky130_fd_sc_hd__nand3_4 _38671_ (.A(_16294_),
    .B(_16290_),
    .C(_16292_),
    .Y(_16306_));
 sky130_fd_sc_hd__nand3_2 _38672_ (.A(_16302_),
    .B(_16305_),
    .C(_16306_),
    .Y(_16307_));
 sky130_fd_sc_hd__nand3_4 _38673_ (.A(_16299_),
    .B(_16301_),
    .C(_16307_),
    .Y(_16308_));
 sky130_fd_sc_hd__o21ai_2 _38674_ (.A1(_16295_),
    .A2(_16298_),
    .B1(_16305_),
    .Y(_16309_));
 sky130_fd_sc_hd__a21boi_2 _38675_ (.A1(_16065_),
    .A2(_16085_),
    .B1_N(_16066_),
    .Y(_16310_));
 sky130_fd_sc_hd__nand3_2 _38676_ (.A(_16302_),
    .B(_16306_),
    .C(_16304_),
    .Y(_16311_));
 sky130_fd_sc_hd__nand3_4 _38677_ (.A(_16309_),
    .B(_16310_),
    .C(_16311_),
    .Y(_16312_));
 sky130_fd_sc_hd__buf_8 _38678_ (.A(_14329_),
    .X(_16313_));
 sky130_fd_sc_hd__nand2_4 _38679_ (.A(_16095_),
    .B(_16078_),
    .Y(_16314_));
 sky130_vsdinv _38680_ (.A(_16314_),
    .Y(_16315_));
 sky130_fd_sc_hd__nor2_8 _38681_ (.A(_16313_),
    .B(_16315_),
    .Y(_16316_));
 sky130_fd_sc_hd__buf_6 _38682_ (.A(_14592_),
    .X(_16317_));
 sky130_fd_sc_hd__buf_6 _38683_ (.A(_16317_),
    .X(_16318_));
 sky130_fd_sc_hd__nor2_1 _38684_ (.A(_16318_),
    .B(_16314_),
    .Y(_16319_));
 sky130_fd_sc_hd__o2bb2ai_2 _38685_ (.A1_N(_16308_),
    .A2_N(_16312_),
    .B1(_16316_),
    .B2(_16319_),
    .Y(_16320_));
 sky130_fd_sc_hd__xor2_4 _38686_ (.A(_16317_),
    .B(_16314_),
    .X(_16321_));
 sky130_fd_sc_hd__nand3_2 _38687_ (.A(_16312_),
    .B(_16308_),
    .C(_16321_),
    .Y(_16322_));
 sky130_fd_sc_hd__nand3_4 _38688_ (.A(_16139_),
    .B(_16320_),
    .C(_16322_),
    .Y(_16323_));
 sky130_fd_sc_hd__nor2_1 _38689_ (.A(_16318_),
    .B(_16315_),
    .Y(_16324_));
 sky130_fd_sc_hd__nor2_1 _38690_ (.A(_14331_),
    .B(_16314_),
    .Y(_16325_));
 sky130_fd_sc_hd__o2bb2ai_2 _38691_ (.A1_N(_16308_),
    .A2_N(_16312_),
    .B1(_16324_),
    .B2(_16325_),
    .Y(_16326_));
 sky130_fd_sc_hd__a21oi_2 _38692_ (.A1(_16098_),
    .A2(_16102_),
    .B1(_16138_),
    .Y(_16327_));
 sky130_fd_sc_hd__nand3b_2 _38693_ (.A_N(_16321_),
    .B(_16312_),
    .C(_16308_),
    .Y(_16328_));
 sky130_fd_sc_hd__nand3_4 _38694_ (.A(_16326_),
    .B(_16327_),
    .C(_16328_),
    .Y(_16329_));
 sky130_fd_sc_hd__buf_2 _38695_ (.A(_16101_),
    .X(_16330_));
 sky130_fd_sc_hd__a21oi_1 _38696_ (.A1(_16323_),
    .A2(_16329_),
    .B1(_16330_),
    .Y(_16331_));
 sky130_fd_sc_hd__and3_1 _38697_ (.A(_16323_),
    .B(_16329_),
    .C(_16330_),
    .X(_16332_));
 sky130_fd_sc_hd__nand2_1 _38698_ (.A(_16108_),
    .B(_16109_),
    .Y(_16333_));
 sky130_fd_sc_hd__a21boi_2 _38699_ (.A1(_16333_),
    .A2(_16105_),
    .B1_N(_15901_),
    .Y(_16334_));
 sky130_fd_sc_hd__nor2_1 _38700_ (.A(_16112_),
    .B(_16334_),
    .Y(_16335_));
 sky130_fd_sc_hd__o21ai_2 _38701_ (.A1(_16331_),
    .A2(_16332_),
    .B1(_16335_),
    .Y(_16336_));
 sky130_fd_sc_hd__nand2_2 _38702_ (.A(_16113_),
    .B(_16110_),
    .Y(_16337_));
 sky130_fd_sc_hd__nand2_1 _38703_ (.A(_16323_),
    .B(_16329_),
    .Y(_16338_));
 sky130_vsdinv _38704_ (.A(_16330_),
    .Y(_16339_));
 sky130_fd_sc_hd__nand2_2 _38705_ (.A(_16338_),
    .B(_16339_),
    .Y(_16340_));
 sky130_fd_sc_hd__nand3_4 _38706_ (.A(_16323_),
    .B(_16329_),
    .C(_16330_),
    .Y(_16341_));
 sky130_fd_sc_hd__nand3_4 _38707_ (.A(_16337_),
    .B(_16340_),
    .C(_16341_),
    .Y(_16342_));
 sky130_fd_sc_hd__and2_2 _38708_ (.A(_16336_),
    .B(_16342_),
    .X(_16343_));
 sky130_fd_sc_hd__nand2_2 _38709_ (.A(_16137_),
    .B(_16118_),
    .Y(_16344_));
 sky130_fd_sc_hd__xor2_4 _38710_ (.A(_16343_),
    .B(_16344_),
    .X(_02668_));
 sky130_fd_sc_hd__o21a_2 _38711_ (.A1(_16304_),
    .A2(_16295_),
    .B1(_16306_),
    .X(_16345_));
 sky130_fd_sc_hd__nand2_1 _38712_ (.A(_16288_),
    .B(_16286_),
    .Y(_16346_));
 sky130_fd_sc_hd__nand3b_4 _38713_ (.A_N(_16286_),
    .B(_16281_),
    .C(_16285_),
    .Y(_16347_));
 sky130_fd_sc_hd__nand2_1 _38714_ (.A(_16346_),
    .B(_16347_),
    .Y(_16348_));
 sky130_fd_sc_hd__nand2_1 _38715_ (.A(_16253_),
    .B(_16348_),
    .Y(_16349_));
 sky130_fd_sc_hd__nor2_4 _38716_ (.A(_15823_),
    .B(_08080_),
    .Y(_16350_));
 sky130_fd_sc_hd__and4_2 _38717_ (.A(_10732_),
    .B(_15937_),
    .C(_19577_),
    .D(_19872_),
    .X(_16351_));
 sky130_fd_sc_hd__clkbuf_2 _38718_ (.A(_13745_),
    .X(_16352_));
 sky130_fd_sc_hd__clkbuf_4 _38719_ (.A(_15939_),
    .X(_16353_));
 sky130_fd_sc_hd__o22a_2 _38720_ (.A1(_19875_),
    .A2(_16352_),
    .B1(_16353_),
    .B2(_10971_),
    .X(_16354_));
 sky130_fd_sc_hd__or3_4 _38721_ (.A(_16350_),
    .B(_16351_),
    .C(_16354_),
    .X(_16355_));
 sky130_fd_sc_hd__o21ai_4 _38722_ (.A1(_16351_),
    .A2(_16354_),
    .B1(_16350_),
    .Y(_16356_));
 sky130_fd_sc_hd__nor2_1 _38723_ (.A(_16169_),
    .B(_16166_),
    .Y(_16357_));
 sky130_fd_sc_hd__or2_4 _38724_ (.A(_16167_),
    .B(_16357_),
    .X(_16358_));
 sky130_fd_sc_hd__a21oi_4 _38725_ (.A1(_16355_),
    .A2(_16356_),
    .B1(_16358_),
    .Y(_16359_));
 sky130_fd_sc_hd__and3_1 _38726_ (.A(_16358_),
    .B(_16355_),
    .C(_16356_),
    .X(_16360_));
 sky130_fd_sc_hd__nand2_4 _38727_ (.A(_15806_),
    .B(_19860_),
    .Y(_16361_));
 sky130_fd_sc_hd__o22a_1 _38728_ (.A1(_16159_),
    .A2(_12916_),
    .B1(_15932_),
    .B2(_12078_),
    .X(_16362_));
 sky130_fd_sc_hd__a31o_2 _38729_ (.A1(_19864_),
    .A2(_19867_),
    .A3(_15930_),
    .B1(_16362_),
    .X(_16363_));
 sky130_fd_sc_hd__nor2_4 _38730_ (.A(_16361_),
    .B(_16363_),
    .Y(_16364_));
 sky130_fd_sc_hd__and2_2 _38731_ (.A(_16363_),
    .B(_16361_),
    .X(_16365_));
 sky130_fd_sc_hd__nor2_8 _38732_ (.A(_16364_),
    .B(_16365_),
    .Y(_16366_));
 sky130_fd_sc_hd__o21ai_2 _38733_ (.A1(_16359_),
    .A2(_16360_),
    .B1(_16366_),
    .Y(_16367_));
 sky130_fd_sc_hd__a21boi_2 _38734_ (.A1(_16165_),
    .A2(_16175_),
    .B1_N(_16176_),
    .Y(_16368_));
 sky130_fd_sc_hd__nand2_1 _38735_ (.A(_16363_),
    .B(_16361_),
    .Y(_16369_));
 sky130_fd_sc_hd__or2b_2 _38736_ (.A(_16364_),
    .B_N(_16369_),
    .X(_16370_));
 sky130_fd_sc_hd__nand3_4 _38737_ (.A(_16358_),
    .B(_16356_),
    .C(_16355_),
    .Y(_16371_));
 sky130_fd_sc_hd__a21o_1 _38738_ (.A1(_16355_),
    .A2(_16356_),
    .B1(_16358_),
    .X(_16372_));
 sky130_fd_sc_hd__nand3_2 _38739_ (.A(_16370_),
    .B(_16371_),
    .C(_16372_),
    .Y(_16373_));
 sky130_fd_sc_hd__nand3_4 _38740_ (.A(_16367_),
    .B(_16368_),
    .C(_16373_),
    .Y(_16374_));
 sky130_fd_sc_hd__o21ai_2 _38741_ (.A1(_16359_),
    .A2(_16360_),
    .B1(_16370_),
    .Y(_16375_));
 sky130_fd_sc_hd__nand2_1 _38742_ (.A(_16177_),
    .B(_16176_),
    .Y(_16376_));
 sky130_fd_sc_hd__nand3_2 _38743_ (.A(_16366_),
    .B(_16372_),
    .C(_16371_),
    .Y(_16377_));
 sky130_fd_sc_hd__nand3_4 _38744_ (.A(_16375_),
    .B(_16376_),
    .C(_16377_),
    .Y(_16378_));
 sky130_fd_sc_hd__or2_2 _38745_ (.A(_16183_),
    .B(_16188_),
    .X(_16379_));
 sky130_fd_sc_hd__nand2_1 _38746_ (.A(_19598_),
    .B(_14501_),
    .Y(_16380_));
 sky130_fd_sc_hd__nand2_1 _38747_ (.A(_19601_),
    .B(_11224_),
    .Y(_16381_));
 sky130_fd_sc_hd__or2_2 _38748_ (.A(_16380_),
    .B(_16381_),
    .X(_16382_));
 sky130_fd_sc_hd__nand2_2 _38749_ (.A(_16380_),
    .B(_16381_),
    .Y(_16383_));
 sky130_fd_sc_hd__nand2_1 _38750_ (.A(_19604_),
    .B(_19850_),
    .Y(_16384_));
 sky130_fd_sc_hd__a21bo_1 _38751_ (.A1(_16382_),
    .A2(_16383_),
    .B1_N(_16384_),
    .X(_16385_));
 sky130_fd_sc_hd__nand3b_4 _38752_ (.A_N(_16384_),
    .B(_16382_),
    .C(_16383_),
    .Y(_16386_));
 sky130_fd_sc_hd__o21bai_4 _38753_ (.A1(_16158_),
    .A2(_16160_),
    .B1_N(_16162_),
    .Y(_16387_));
 sky130_fd_sc_hd__a21oi_4 _38754_ (.A1(_16385_),
    .A2(_16386_),
    .B1(_16387_),
    .Y(_16388_));
 sky130_fd_sc_hd__and3_2 _38755_ (.A(_16387_),
    .B(_16385_),
    .C(_16386_),
    .X(_16389_));
 sky130_fd_sc_hd__nor2_1 _38756_ (.A(_16388_),
    .B(_16389_),
    .Y(_16390_));
 sky130_fd_sc_hd__nor2_2 _38757_ (.A(_16379_),
    .B(_16390_),
    .Y(_16391_));
 sky130_fd_sc_hd__and2_1 _38758_ (.A(_16390_),
    .B(_16379_),
    .X(_16392_));
 sky130_fd_sc_hd__o2bb2ai_4 _38759_ (.A1_N(_16374_),
    .A2_N(_16378_),
    .B1(_16391_),
    .B2(_16392_),
    .Y(_16393_));
 sky130_fd_sc_hd__nor3_4 _38760_ (.A(_16388_),
    .B(_16379_),
    .C(_16389_),
    .Y(_16394_));
 sky130_fd_sc_hd__o21ai_1 _38761_ (.A1(_16388_),
    .A2(_16389_),
    .B1(_16379_),
    .Y(_16395_));
 sky130_fd_sc_hd__or2b_2 _38762_ (.A(_16394_),
    .B_N(_16395_),
    .X(_16396_));
 sky130_fd_sc_hd__nand3_4 _38763_ (.A(_16396_),
    .B(_16378_),
    .C(_16374_),
    .Y(_16397_));
 sky130_fd_sc_hd__a21oi_4 _38764_ (.A1(_16179_),
    .A2(_16177_),
    .B1(_16157_),
    .Y(_16398_));
 sky130_fd_sc_hd__o21ai_4 _38765_ (.A1(_16205_),
    .A2(_16398_),
    .B1(_16180_),
    .Y(_16399_));
 sky130_fd_sc_hd__a21oi_4 _38766_ (.A1(_16393_),
    .A2(_16397_),
    .B1(_16399_),
    .Y(_16400_));
 sky130_fd_sc_hd__and3_2 _38767_ (.A(_16399_),
    .B(_16393_),
    .C(_16397_),
    .X(_16401_));
 sky130_fd_sc_hd__nand2_1 _38768_ (.A(_19618_),
    .B(_11582_),
    .Y(_16402_));
 sky130_fd_sc_hd__nand2_1 _38769_ (.A(_15769_),
    .B(_10493_),
    .Y(_16403_));
 sky130_fd_sc_hd__nand2_1 _38770_ (.A(_15768_),
    .B(_11574_),
    .Y(_16404_));
 sky130_fd_sc_hd__nor2_2 _38771_ (.A(_16403_),
    .B(_16404_),
    .Y(_16405_));
 sky130_fd_sc_hd__nand2_1 _38772_ (.A(_16403_),
    .B(_16404_),
    .Y(_16406_));
 sky130_fd_sc_hd__or3b_4 _38773_ (.A(_16402_),
    .B(_16405_),
    .C_N(_16406_),
    .X(_16407_));
 sky130_vsdinv _38774_ (.A(_16405_),
    .Y(_16408_));
 sky130_fd_sc_hd__a21bo_1 _38775_ (.A1(_16408_),
    .A2(_16406_),
    .B1_N(_16402_),
    .X(_16409_));
 sky130_fd_sc_hd__nand2_2 _38776_ (.A(_16220_),
    .B(_16216_),
    .Y(_16410_));
 sky130_fd_sc_hd__a21o_1 _38777_ (.A1(_16407_),
    .A2(_16409_),
    .B1(_16410_),
    .X(_16411_));
 sky130_fd_sc_hd__nand3_4 _38778_ (.A(_16407_),
    .B(_16409_),
    .C(_16410_),
    .Y(_16412_));
 sky130_fd_sc_hd__nor2_8 _38779_ (.A(_18468_),
    .B(_07041_),
    .Y(_16413_));
 sky130_fd_sc_hd__and4_4 _38780_ (.A(_11847_),
    .B(_11849_),
    .C(_19825_),
    .D(_11202_),
    .X(_16414_));
 sky130_fd_sc_hd__o21a_1 _38781_ (.A1(_15993_),
    .A2(_12618_),
    .B1(_16225_),
    .X(_16415_));
 sky130_fd_sc_hd__nor2_1 _38782_ (.A(_16414_),
    .B(_16415_),
    .Y(_16416_));
 sky130_fd_sc_hd__nor2_1 _38783_ (.A(_16413_),
    .B(_16416_),
    .Y(_16417_));
 sky130_fd_sc_hd__and2_1 _38784_ (.A(_16416_),
    .B(_16413_),
    .X(_16418_));
 sky130_fd_sc_hd__nor2_2 _38785_ (.A(_16417_),
    .B(_16418_),
    .Y(_16419_));
 sky130_fd_sc_hd__a21o_1 _38786_ (.A1(_16411_),
    .A2(_16412_),
    .B1(_16419_),
    .X(_16420_));
 sky130_fd_sc_hd__nand3_4 _38787_ (.A(_16411_),
    .B(_16412_),
    .C(_16419_),
    .Y(_16421_));
 sky130_fd_sc_hd__o21ai_2 _38788_ (.A1(_16196_),
    .A2(_16192_),
    .B1(_16199_),
    .Y(_16422_));
 sky130_fd_sc_hd__a21o_2 _38789_ (.A1(_16420_),
    .A2(_16421_),
    .B1(_16422_),
    .X(_16423_));
 sky130_fd_sc_hd__nand3_4 _38790_ (.A(_16422_),
    .B(_16420_),
    .C(_16421_),
    .Y(_16424_));
 sky130_fd_sc_hd__nand2_4 _38791_ (.A(_16233_),
    .B(_16223_),
    .Y(_16425_));
 sky130_fd_sc_hd__a21o_1 _38792_ (.A1(_16423_),
    .A2(_16424_),
    .B1(_16425_),
    .X(_16426_));
 sky130_fd_sc_hd__nand3_4 _38793_ (.A(_16423_),
    .B(_16424_),
    .C(_16425_),
    .Y(_16427_));
 sky130_fd_sc_hd__nand2_4 _38794_ (.A(_16426_),
    .B(_16427_),
    .Y(_16428_));
 sky130_fd_sc_hd__o21ai_4 _38795_ (.A1(_16400_),
    .A2(_16401_),
    .B1(_16428_),
    .Y(_16429_));
 sky130_fd_sc_hd__o21ai_4 _38796_ (.A1(_16246_),
    .A2(_16208_),
    .B1(_16245_),
    .Y(_16430_));
 sky130_fd_sc_hd__a21o_2 _38797_ (.A1(_16393_),
    .A2(_16397_),
    .B1(_16399_),
    .X(_16431_));
 sky130_fd_sc_hd__a21oi_4 _38798_ (.A1(_16423_),
    .A2(_16424_),
    .B1(_16425_),
    .Y(_16432_));
 sky130_fd_sc_hd__and3_2 _38799_ (.A(_16423_),
    .B(_16424_),
    .C(_16425_),
    .X(_16433_));
 sky130_fd_sc_hd__nor2_8 _38800_ (.A(_16432_),
    .B(_16433_),
    .Y(_16434_));
 sky130_fd_sc_hd__nand3_4 _38801_ (.A(_16399_),
    .B(_16393_),
    .C(_16397_),
    .Y(_16435_));
 sky130_fd_sc_hd__nand3_4 _38802_ (.A(_16431_),
    .B(_16434_),
    .C(_16435_),
    .Y(_16436_));
 sky130_fd_sc_hd__nand3_4 _38803_ (.A(_16429_),
    .B(_16430_),
    .C(_16436_),
    .Y(_16437_));
 sky130_fd_sc_hd__o21ai_2 _38804_ (.A1(_16400_),
    .A2(_16401_),
    .B1(_16434_),
    .Y(_16438_));
 sky130_fd_sc_hd__a21oi_4 _38805_ (.A1(_16244_),
    .A2(_16241_),
    .B1(_16211_),
    .Y(_16439_));
 sky130_fd_sc_hd__nand3_4 _38806_ (.A(_16431_),
    .B(_16435_),
    .C(_16428_),
    .Y(_16440_));
 sky130_fd_sc_hd__nand3_4 _38807_ (.A(_16438_),
    .B(_16439_),
    .C(_16440_),
    .Y(_16441_));
 sky130_fd_sc_hd__nor2_4 _38808_ (.A(_16266_),
    .B(_16265_),
    .Y(_16442_));
 sky130_fd_sc_hd__nor2_4 _38809_ (.A(_15995_),
    .B(_16225_),
    .Y(_16443_));
 sky130_fd_sc_hd__o21ai_4 _38810_ (.A1(_16443_),
    .A2(_16229_),
    .B1(_16265_),
    .Y(_16444_));
 sky130_fd_sc_hd__a211o_2 _38811_ (.A1(_16260_),
    .A2(_16262_),
    .B1(_16443_),
    .C1(_16229_),
    .X(_16445_));
 sky130_vsdinv _38812_ (.A(_16257_),
    .Y(_16446_));
 sky130_fd_sc_hd__nand2_4 _38813_ (.A(_16446_),
    .B(_16259_),
    .Y(_16447_));
 sky130_vsdinv _38814_ (.A(_16447_),
    .Y(_16448_));
 sky130_fd_sc_hd__nand3_2 _38815_ (.A(_16444_),
    .B(_16445_),
    .C(_16448_),
    .Y(_16449_));
 sky130_fd_sc_hd__nand2_1 _38816_ (.A(_16444_),
    .B(_16445_),
    .Y(_16450_));
 sky130_fd_sc_hd__nand2_1 _38817_ (.A(_16450_),
    .B(_16447_),
    .Y(_16451_));
 sky130_fd_sc_hd__o2111ai_4 _38818_ (.A1(_16270_),
    .A2(_16442_),
    .B1(_16267_),
    .C1(_16449_),
    .D1(_16451_),
    .Y(_16452_));
 sky130_fd_sc_hd__nand2_1 _38819_ (.A(_16450_),
    .B(_16448_),
    .Y(_16453_));
 sky130_fd_sc_hd__o21ai_2 _38820_ (.A1(_16270_),
    .A2(_16442_),
    .B1(_16267_),
    .Y(_16454_));
 sky130_fd_sc_hd__nand3_2 _38821_ (.A(_16444_),
    .B(_16445_),
    .C(_16447_),
    .Y(_16455_));
 sky130_fd_sc_hd__nand3_4 _38822_ (.A(_16453_),
    .B(_16454_),
    .C(_16455_),
    .Y(_16456_));
 sky130_fd_sc_hd__nand3_2 _38823_ (.A(_16452_),
    .B(_16456_),
    .C(_16045_),
    .Y(_16457_));
 sky130_fd_sc_hd__nand2_1 _38824_ (.A(_16452_),
    .B(_16456_),
    .Y(_16458_));
 sky130_fd_sc_hd__nand2_1 _38825_ (.A(_16458_),
    .B(_16048_),
    .Y(_16459_));
 sky130_fd_sc_hd__o2111ai_4 _38826_ (.A1(_16235_),
    .A2(_16236_),
    .B1(_16457_),
    .C1(_16240_),
    .D1(_16459_),
    .Y(_16460_));
 sky130_fd_sc_hd__nand2_1 _38827_ (.A(_16240_),
    .B(_16234_),
    .Y(_16461_));
 sky130_fd_sc_hd__nand2_1 _38828_ (.A(_16458_),
    .B(_16045_),
    .Y(_16462_));
 sky130_fd_sc_hd__nand3_2 _38829_ (.A(_16452_),
    .B(_16456_),
    .C(_16048_),
    .Y(_16463_));
 sky130_fd_sc_hd__nand3_4 _38830_ (.A(_16461_),
    .B(_16462_),
    .C(_16463_),
    .Y(_16464_));
 sky130_fd_sc_hd__nand2_1 _38831_ (.A(_16274_),
    .B(_16048_),
    .Y(_16465_));
 sky130_fd_sc_hd__nand2_2 _38832_ (.A(_16465_),
    .B(_16277_),
    .Y(_16466_));
 sky130_fd_sc_hd__a21o_1 _38833_ (.A1(_16460_),
    .A2(_16464_),
    .B1(_16466_),
    .X(_16467_));
 sky130_vsdinv _38834_ (.A(_16467_),
    .Y(_16468_));
 sky130_fd_sc_hd__nand3_4 _38835_ (.A(_16460_),
    .B(_16464_),
    .C(_16466_),
    .Y(_16469_));
 sky130_vsdinv _38836_ (.A(_16469_),
    .Y(_16470_));
 sky130_fd_sc_hd__o2bb2ai_4 _38837_ (.A1_N(_16437_),
    .A2_N(_16441_),
    .B1(_16468_),
    .B2(_16470_),
    .Y(_16471_));
 sky130_fd_sc_hd__nand2_2 _38838_ (.A(_16467_),
    .B(_16469_),
    .Y(_16472_));
 sky130_fd_sc_hd__nand3b_4 _38839_ (.A_N(_16472_),
    .B(_16441_),
    .C(_16437_),
    .Y(_16473_));
 sky130_fd_sc_hd__a22oi_4 _38840_ (.A1(_16248_),
    .A2(_16349_),
    .B1(_16471_),
    .B2(_16473_),
    .Y(_16474_));
 sky130_fd_sc_hd__a31oi_1 _38841_ (.A1(_16242_),
    .A2(_16247_),
    .A3(_16243_),
    .B1(_16348_),
    .Y(_16475_));
 sky130_fd_sc_hd__o211a_1 _38842_ (.A1(_16296_),
    .A2(_16475_),
    .B1(_16473_),
    .C1(_16471_),
    .X(_16476_));
 sky130_fd_sc_hd__a21o_1 _38843_ (.A1(_16347_),
    .A2(_16285_),
    .B1(_16149_),
    .X(_16477_));
 sky130_fd_sc_hd__buf_4 _38844_ (.A(_16148_),
    .X(_16478_));
 sky130_fd_sc_hd__nand3_4 _38845_ (.A(_16347_),
    .B(_16478_),
    .C(_16285_),
    .Y(_16479_));
 sky130_fd_sc_hd__nor2_4 _38846_ (.A(_16141_),
    .B(_13989_),
    .Y(_16480_));
 sky130_fd_sc_hd__nor2_1 _38847_ (.A(_16145_),
    .B(_16480_),
    .Y(_16481_));
 sky130_fd_sc_hd__buf_2 _38848_ (.A(_16481_),
    .X(_16482_));
 sky130_fd_sc_hd__a21o_1 _38849_ (.A1(_16477_),
    .A2(_16479_),
    .B1(_16482_),
    .X(_16483_));
 sky130_fd_sc_hd__buf_4 _38850_ (.A(_16481_),
    .X(_16484_));
 sky130_fd_sc_hd__nand3_4 _38851_ (.A(_16477_),
    .B(_16479_),
    .C(_16484_),
    .Y(_16485_));
 sky130_fd_sc_hd__and2_2 _38852_ (.A(_16483_),
    .B(_16485_),
    .X(_16486_));
 sky130_fd_sc_hd__o21ai_4 _38853_ (.A1(_16474_),
    .A2(_16476_),
    .B1(_16486_),
    .Y(_16487_));
 sky130_fd_sc_hd__nand2_2 _38854_ (.A(_16297_),
    .B(_16253_),
    .Y(_16488_));
 sky130_fd_sc_hd__a21o_2 _38855_ (.A1(_16471_),
    .A2(_16473_),
    .B1(_16488_),
    .X(_16489_));
 sky130_fd_sc_hd__nand2_4 _38856_ (.A(_16483_),
    .B(_16485_),
    .Y(_16490_));
 sky130_fd_sc_hd__nand3_4 _38857_ (.A(_16488_),
    .B(_16471_),
    .C(_16473_),
    .Y(_16491_));
 sky130_fd_sc_hd__nand3_4 _38858_ (.A(_16489_),
    .B(_16490_),
    .C(_16491_),
    .Y(_16492_));
 sky130_fd_sc_hd__nand3_4 _38859_ (.A(_16345_),
    .B(_16487_),
    .C(_16492_),
    .Y(_16493_));
 sky130_fd_sc_hd__o21ai_2 _38860_ (.A1(_16474_),
    .A2(_16476_),
    .B1(_16490_),
    .Y(_16494_));
 sky130_fd_sc_hd__o21ai_2 _38861_ (.A1(_16304_),
    .A2(_16295_),
    .B1(_16306_),
    .Y(_16495_));
 sky130_fd_sc_hd__nand3_4 _38862_ (.A(_16489_),
    .B(_16486_),
    .C(_16491_),
    .Y(_16496_));
 sky130_fd_sc_hd__nand3_4 _38863_ (.A(_16494_),
    .B(_16495_),
    .C(_16496_),
    .Y(_16497_));
 sky130_fd_sc_hd__nand2_2 _38864_ (.A(_16155_),
    .B(_16150_),
    .Y(_16498_));
 sky130_fd_sc_hd__nor2_4 _38865_ (.A(_14330_),
    .B(_16498_),
    .Y(_16499_));
 sky130_vsdinv _38866_ (.A(_16498_),
    .Y(_16500_));
 sky130_fd_sc_hd__nor2_4 _38867_ (.A(_16317_),
    .B(_16500_),
    .Y(_16501_));
 sky130_fd_sc_hd__or2_2 _38868_ (.A(_16499_),
    .B(_16501_),
    .X(_16502_));
 sky130_fd_sc_hd__a21o_1 _38869_ (.A1(_16493_),
    .A2(_16497_),
    .B1(_16502_),
    .X(_16503_));
 sky130_fd_sc_hd__nand2_1 _38870_ (.A(_16312_),
    .B(_16321_),
    .Y(_16504_));
 sky130_fd_sc_hd__nand2_1 _38871_ (.A(_16504_),
    .B(_16308_),
    .Y(_16505_));
 sky130_fd_sc_hd__nand3_2 _38872_ (.A(_16493_),
    .B(_16497_),
    .C(_16502_),
    .Y(_16506_));
 sky130_fd_sc_hd__nand3_4 _38873_ (.A(_16503_),
    .B(_16505_),
    .C(_16506_),
    .Y(_16507_));
 sky130_fd_sc_hd__o2bb2ai_4 _38874_ (.A1_N(_16497_),
    .A2_N(_16493_),
    .B1(_16501_),
    .B2(_16499_),
    .Y(_16508_));
 sky130_fd_sc_hd__a21boi_4 _38875_ (.A1(_16312_),
    .A2(_16321_),
    .B1_N(_16308_),
    .Y(_16509_));
 sky130_fd_sc_hd__nor2_4 _38876_ (.A(_16499_),
    .B(_16501_),
    .Y(_16510_));
 sky130_fd_sc_hd__nand3_4 _38877_ (.A(_16493_),
    .B(_16497_),
    .C(_16510_),
    .Y(_16511_));
 sky130_fd_sc_hd__nand3_4 _38878_ (.A(_16508_),
    .B(_16509_),
    .C(_16511_),
    .Y(_16512_));
 sky130_fd_sc_hd__nand3_4 _38879_ (.A(_16507_),
    .B(_16512_),
    .C(_16316_),
    .Y(_16513_));
 sky130_vsdinv _38880_ (.A(_16513_),
    .Y(_16514_));
 sky130_fd_sc_hd__buf_6 _38881_ (.A(net410),
    .X(_16515_));
 sky130_fd_sc_hd__o2bb2ai_2 _38882_ (.A1_N(_16512_),
    .A2_N(_16507_),
    .B1(_16515_),
    .B2(_16315_),
    .Y(_16516_));
 sky130_fd_sc_hd__nand2_1 _38883_ (.A(_16329_),
    .B(_16330_),
    .Y(_16517_));
 sky130_fd_sc_hd__nand2_2 _38884_ (.A(_16517_),
    .B(_16323_),
    .Y(_16518_));
 sky130_fd_sc_hd__nand2_1 _38885_ (.A(_16516_),
    .B(_16518_),
    .Y(_16519_));
 sky130_vsdinv _38886_ (.A(_16316_),
    .Y(_16520_));
 sky130_fd_sc_hd__a21o_1 _38887_ (.A1(_16507_),
    .A2(_16512_),
    .B1(_16520_),
    .X(_16521_));
 sky130_fd_sc_hd__a21boi_2 _38888_ (.A1(_16330_),
    .A2(_16329_),
    .B1_N(_16323_),
    .Y(_16522_));
 sky130_fd_sc_hd__nand3_2 _38889_ (.A(_16507_),
    .B(_16512_),
    .C(_16520_),
    .Y(_16523_));
 sky130_fd_sc_hd__nand3_4 _38890_ (.A(_16521_),
    .B(_16522_),
    .C(_16523_),
    .Y(_16524_));
 sky130_fd_sc_hd__o21a_2 _38891_ (.A1(_16514_),
    .A2(_16519_),
    .B1(_16524_),
    .X(_16525_));
 sky130_fd_sc_hd__o2bb2ai_2 _38892_ (.A1_N(_16339_),
    .A2_N(_16338_),
    .B1(_16112_),
    .B2(_16334_),
    .Y(_16526_));
 sky130_fd_sc_hd__o2111ai_4 _38893_ (.A1(_16332_),
    .A2(_16526_),
    .B1(_16118_),
    .C1(_16336_),
    .D1(_16116_),
    .Y(_16527_));
 sky130_vsdinv _38894_ (.A(_16527_),
    .Y(_16528_));
 sky130_fd_sc_hd__a21oi_2 _38895_ (.A1(_16340_),
    .A2(_16341_),
    .B1(_16337_),
    .Y(_16529_));
 sky130_fd_sc_hd__a21oi_4 _38896_ (.A1(_16118_),
    .A2(_16342_),
    .B1(_16529_),
    .Y(_16530_));
 sky130_fd_sc_hd__a21oi_4 _38897_ (.A1(_16135_),
    .A2(_16528_),
    .B1(_16530_),
    .Y(_16531_));
 sky130_fd_sc_hd__xnor2_4 _38898_ (.A(_16525_),
    .B(_16531_),
    .Y(_02669_));
 sky130_fd_sc_hd__and3_1 _38899_ (.A(_16494_),
    .B(_16496_),
    .C(_16495_),
    .X(_16532_));
 sky130_fd_sc_hd__a31oi_4 _38900_ (.A1(_16345_),
    .A2(_16487_),
    .A3(_16492_),
    .B1(_16510_),
    .Y(_16533_));
 sky130_fd_sc_hd__nor2_4 _38901_ (.A(_15823_),
    .B(_12916_),
    .Y(_16534_));
 sky130_fd_sc_hd__and4_2 _38902_ (.A(_11694_),
    .B(_15937_),
    .C(_15821_),
    .D(_11724_),
    .X(_16535_));
 sky130_fd_sc_hd__o22a_2 _38903_ (.A1(_19872_),
    .A2(_16352_),
    .B1(_15817_),
    .B2(_08080_),
    .X(_16536_));
 sky130_fd_sc_hd__or3_4 _38904_ (.A(_16534_),
    .B(_16535_),
    .C(_16536_),
    .X(_16537_));
 sky130_fd_sc_hd__o21ai_4 _38905_ (.A1(_16535_),
    .A2(_16536_),
    .B1(_16534_),
    .Y(_16538_));
 sky130_fd_sc_hd__nor2_1 _38906_ (.A(_16350_),
    .B(_16351_),
    .Y(_16539_));
 sky130_fd_sc_hd__or2_4 _38907_ (.A(_16354_),
    .B(_16539_),
    .X(_16540_));
 sky130_fd_sc_hd__a21oi_4 _38908_ (.A1(_16537_),
    .A2(_16538_),
    .B1(_16540_),
    .Y(_16541_));
 sky130_fd_sc_hd__o22a_2 _38909_ (.A1(_15931_),
    .A2(net439),
    .B1(_15932_),
    .B2(_10466_),
    .X(_16542_));
 sky130_fd_sc_hd__a31o_1 _38910_ (.A1(_19860_),
    .A2(_19864_),
    .A3(_15930_),
    .B1(_16542_),
    .X(_16543_));
 sky130_fd_sc_hd__nand2_2 _38911_ (.A(_19593_),
    .B(_19856_),
    .Y(_16544_));
 sky130_fd_sc_hd__nand2_2 _38912_ (.A(_16543_),
    .B(_16544_),
    .Y(_16545_));
 sky130_fd_sc_hd__and3_1 _38913_ (.A(_15929_),
    .B(_19859_),
    .C(_10981_),
    .X(_16546_));
 sky130_fd_sc_hd__nor2_1 _38914_ (.A(_16542_),
    .B(_16546_),
    .Y(_16547_));
 sky130_vsdinv _38915_ (.A(_16544_),
    .Y(_16548_));
 sky130_fd_sc_hd__nand2_2 _38916_ (.A(_16547_),
    .B(_16548_),
    .Y(_16549_));
 sky130_fd_sc_hd__and2_1 _38917_ (.A(_16545_),
    .B(_16549_),
    .X(_16550_));
 sky130_fd_sc_hd__nand3_4 _38918_ (.A(_16540_),
    .B(_16538_),
    .C(_16537_),
    .Y(_16551_));
 sky130_fd_sc_hd__nand2_2 _38919_ (.A(_16550_),
    .B(_16551_),
    .Y(_16552_));
 sky130_fd_sc_hd__and3_1 _38920_ (.A(_16540_),
    .B(_16537_),
    .C(_16538_),
    .X(_16553_));
 sky130_fd_sc_hd__nand2_2 _38921_ (.A(_16545_),
    .B(_16549_),
    .Y(_16554_));
 sky130_fd_sc_hd__o21ai_2 _38922_ (.A1(_16541_),
    .A2(_16553_),
    .B1(_16554_),
    .Y(_16555_));
 sky130_fd_sc_hd__a21o_1 _38923_ (.A1(_16366_),
    .A2(_16371_),
    .B1(_16359_),
    .X(_16556_));
 sky130_fd_sc_hd__o211ai_4 _38924_ (.A1(_16541_),
    .A2(_16552_),
    .B1(_16555_),
    .C1(_16556_),
    .Y(_16557_));
 sky130_fd_sc_hd__o21ai_4 _38925_ (.A1(_16541_),
    .A2(_16553_),
    .B1(_16550_),
    .Y(_16558_));
 sky130_fd_sc_hd__a21oi_4 _38926_ (.A1(_16366_),
    .A2(_16371_),
    .B1(_16359_),
    .Y(_16559_));
 sky130_fd_sc_hd__a21o_2 _38927_ (.A1(_16537_),
    .A2(_16538_),
    .B1(_16540_),
    .X(_16560_));
 sky130_fd_sc_hd__nand3_4 _38928_ (.A(_16560_),
    .B(_16551_),
    .C(_16554_),
    .Y(_16561_));
 sky130_fd_sc_hd__nand3_4 _38929_ (.A(_16558_),
    .B(_16559_),
    .C(_16561_),
    .Y(_16562_));
 sky130_fd_sc_hd__and4_2 _38930_ (.A(_13514_),
    .B(_08947_),
    .C(_09359_),
    .D(_09362_),
    .X(_16563_));
 sky130_fd_sc_hd__nand2_2 _38931_ (.A(_13514_),
    .B(_09823_),
    .Y(_16564_));
 sky130_fd_sc_hd__o21a_1 _38932_ (.A1(_15957_),
    .A2(_10617_),
    .B1(_16564_),
    .X(_16565_));
 sky130_fd_sc_hd__nor2_2 _38933_ (.A(_16563_),
    .B(_16565_),
    .Y(_16566_));
 sky130_fd_sc_hd__nand3_4 _38934_ (.A(_16566_),
    .B(_19604_),
    .C(_19845_),
    .Y(_16567_));
 sky130_fd_sc_hd__o32ai_4 _38935_ (.A1(_12078_),
    .A2(_12916_),
    .A3(_15928_),
    .B1(_16361_),
    .B2(_16362_),
    .Y(_16568_));
 sky130_fd_sc_hd__and2_1 _38936_ (.A(_16567_),
    .B(_16568_),
    .X(_16569_));
 sky130_fd_sc_hd__a21o_1 _38937_ (.A1(_19605_),
    .A2(_19846_),
    .B1(_16566_),
    .X(_16570_));
 sky130_fd_sc_hd__nand2_2 _38938_ (.A(_16386_),
    .B(_16382_),
    .Y(_16571_));
 sky130_fd_sc_hd__a21oi_4 _38939_ (.A1(_16570_),
    .A2(_16567_),
    .B1(_16568_),
    .Y(_16572_));
 sky130_fd_sc_hd__a211o_1 _38940_ (.A1(_16569_),
    .A2(_16570_),
    .B1(_16571_),
    .C1(_16572_),
    .X(_16573_));
 sky130_fd_sc_hd__nand3_2 _38941_ (.A(_16570_),
    .B(_16568_),
    .C(_16567_),
    .Y(_16574_));
 sky130_vsdinv _38942_ (.A(_16574_),
    .Y(_16575_));
 sky130_fd_sc_hd__o21ai_2 _38943_ (.A1(_16572_),
    .A2(_16575_),
    .B1(_16571_),
    .Y(_16576_));
 sky130_fd_sc_hd__nand2_4 _38944_ (.A(_16573_),
    .B(_16576_),
    .Y(_16577_));
 sky130_fd_sc_hd__a21o_2 _38945_ (.A1(_16557_),
    .A2(_16562_),
    .B1(_16577_),
    .X(_16578_));
 sky130_fd_sc_hd__nand3_4 _38946_ (.A(_16557_),
    .B(_16577_),
    .C(_16562_),
    .Y(_16579_));
 sky130_fd_sc_hd__nand2_1 _38947_ (.A(_16396_),
    .B(_16374_),
    .Y(_16580_));
 sky130_fd_sc_hd__nand2_4 _38948_ (.A(_16580_),
    .B(_16378_),
    .Y(_16581_));
 sky130_fd_sc_hd__a21oi_4 _38949_ (.A1(_16578_),
    .A2(_16579_),
    .B1(_16581_),
    .Y(_16582_));
 sky130_vsdinv _38950_ (.A(_16378_),
    .Y(_16583_));
 sky130_vsdinv _38951_ (.A(_16395_),
    .Y(_16584_));
 sky130_fd_sc_hd__o21a_1 _38952_ (.A1(_16394_),
    .A2(_16584_),
    .B1(_16374_),
    .X(_16585_));
 sky130_fd_sc_hd__o211a_1 _38953_ (.A1(_16583_),
    .A2(_16585_),
    .B1(_16579_),
    .C1(_16578_),
    .X(_16586_));
 sky130_fd_sc_hd__nand2_2 _38954_ (.A(_19619_),
    .B(_19831_),
    .Y(_16587_));
 sky130_fd_sc_hd__nand2_1 _38955_ (.A(_15769_),
    .B(_19840_),
    .Y(_16588_));
 sky130_fd_sc_hd__nand2_1 _38956_ (.A(_15768_),
    .B(_19835_),
    .Y(_16589_));
 sky130_fd_sc_hd__nor2_2 _38957_ (.A(_16588_),
    .B(_16589_),
    .Y(_16590_));
 sky130_fd_sc_hd__and2_1 _38958_ (.A(_16588_),
    .B(_16589_),
    .X(_16591_));
 sky130_fd_sc_hd__or3_4 _38959_ (.A(_16587_),
    .B(_16590_),
    .C(_16591_),
    .X(_16592_));
 sky130_fd_sc_hd__o21ai_2 _38960_ (.A1(_16590_),
    .A2(_16591_),
    .B1(_16587_),
    .Y(_16593_));
 sky130_fd_sc_hd__a31oi_2 _38961_ (.A1(_16406_),
    .A2(_19619_),
    .A3(_19837_),
    .B1(_16405_),
    .Y(_16594_));
 sky130_fd_sc_hd__a21bo_1 _38962_ (.A1(_16592_),
    .A2(_16593_),
    .B1_N(_16594_),
    .X(_16595_));
 sky130_fd_sc_hd__nand3b_4 _38963_ (.A_N(_16594_),
    .B(_16592_),
    .C(_16593_),
    .Y(_16596_));
 sky130_fd_sc_hd__and4_2 _38964_ (.A(_11594_),
    .B(_19623_),
    .C(_19626_),
    .D(_19826_),
    .X(_16597_));
 sky130_fd_sc_hd__nand2_2 _38965_ (.A(_11593_),
    .B(_19625_),
    .Y(_16598_));
 sky130_fd_sc_hd__o21a_2 _38966_ (.A1(_15992_),
    .A2(_13007_),
    .B1(_16598_),
    .X(_16599_));
 sky130_fd_sc_hd__nor2_4 _38967_ (.A(_16597_),
    .B(_16599_),
    .Y(_16600_));
 sky130_fd_sc_hd__xor2_4 _38968_ (.A(_16413_),
    .B(_16600_),
    .X(_16601_));
 sky130_fd_sc_hd__a21o_1 _38969_ (.A1(_16595_),
    .A2(_16596_),
    .B1(_16601_),
    .X(_16602_));
 sky130_fd_sc_hd__nand3_4 _38970_ (.A(_16595_),
    .B(_16601_),
    .C(_16596_),
    .Y(_16603_));
 sky130_fd_sc_hd__nor2_2 _38971_ (.A(_16183_),
    .B(_16188_),
    .Y(_16604_));
 sky130_fd_sc_hd__o21bai_4 _38972_ (.A1(_16604_),
    .A2(_16388_),
    .B1_N(_16389_),
    .Y(_16605_));
 sky130_fd_sc_hd__a21o_1 _38973_ (.A1(_16602_),
    .A2(_16603_),
    .B1(_16605_),
    .X(_16606_));
 sky130_fd_sc_hd__nand3_4 _38974_ (.A(_16602_),
    .B(_16605_),
    .C(_16603_),
    .Y(_16607_));
 sky130_fd_sc_hd__nand2_1 _38975_ (.A(_16421_),
    .B(_16412_),
    .Y(_16608_));
 sky130_fd_sc_hd__and2_1 _38976_ (.A(_16607_),
    .B(_16608_),
    .X(_16609_));
 sky130_fd_sc_hd__a21oi_2 _38977_ (.A1(_16606_),
    .A2(_16607_),
    .B1(_16608_),
    .Y(_16610_));
 sky130_fd_sc_hd__a21o_2 _38978_ (.A1(_16606_),
    .A2(_16609_),
    .B1(_16610_),
    .X(_16611_));
 sky130_fd_sc_hd__o21ai_2 _38979_ (.A1(_16582_),
    .A2(_16586_),
    .B1(_16611_),
    .Y(_16612_));
 sky130_fd_sc_hd__o21ai_2 _38980_ (.A1(_16428_),
    .A2(_16400_),
    .B1(_16435_),
    .Y(_16613_));
 sky130_fd_sc_hd__a21o_1 _38981_ (.A1(_16578_),
    .A2(_16579_),
    .B1(_16581_),
    .X(_16614_));
 sky130_fd_sc_hd__nand3_4 _38982_ (.A(_16581_),
    .B(_16578_),
    .C(_16579_),
    .Y(_16615_));
 sky130_fd_sc_hd__a21oi_2 _38983_ (.A1(_16606_),
    .A2(_16609_),
    .B1(_16610_),
    .Y(_16616_));
 sky130_fd_sc_hd__nand3_2 _38984_ (.A(_16614_),
    .B(_16615_),
    .C(_16616_),
    .Y(_16617_));
 sky130_fd_sc_hd__nand3_4 _38985_ (.A(_16612_),
    .B(_16613_),
    .C(_16617_),
    .Y(_16618_));
 sky130_fd_sc_hd__o21ai_2 _38986_ (.A1(_16582_),
    .A2(_16586_),
    .B1(_16616_),
    .Y(_16619_));
 sky130_fd_sc_hd__a21oi_4 _38987_ (.A1(_16431_),
    .A2(_16434_),
    .B1(_16401_),
    .Y(_16620_));
 sky130_fd_sc_hd__nand3_4 _38988_ (.A(_16614_),
    .B(_16615_),
    .C(_16611_),
    .Y(_16621_));
 sky130_fd_sc_hd__nand3_4 _38989_ (.A(_16619_),
    .B(_16620_),
    .C(_16621_),
    .Y(_16622_));
 sky130_fd_sc_hd__o21ai_4 _38990_ (.A1(_16414_),
    .A2(_16418_),
    .B1(_16265_),
    .Y(_16623_));
 sky130_fd_sc_hd__nand2_1 _38991_ (.A(_16416_),
    .B(_16413_),
    .Y(_16624_));
 sky130_fd_sc_hd__nand3b_4 _38992_ (.A_N(_16414_),
    .B(_16263_),
    .C(_16624_),
    .Y(_16625_));
 sky130_fd_sc_hd__a21o_1 _38993_ (.A1(_16623_),
    .A2(_16625_),
    .B1(_16447_),
    .X(_16626_));
 sky130_fd_sc_hd__nand3_4 _38994_ (.A(_16623_),
    .B(_16625_),
    .C(_16447_),
    .Y(_16627_));
 sky130_fd_sc_hd__nand2_1 _38995_ (.A(_16445_),
    .B(_16447_),
    .Y(_16628_));
 sky130_fd_sc_hd__nand2_2 _38996_ (.A(_16628_),
    .B(_16444_),
    .Y(_16629_));
 sky130_fd_sc_hd__a21oi_4 _38997_ (.A1(_16626_),
    .A2(_16627_),
    .B1(_16629_),
    .Y(_16630_));
 sky130_fd_sc_hd__nand3_2 _38998_ (.A(_16626_),
    .B(_16629_),
    .C(_16627_),
    .Y(_16631_));
 sky130_fd_sc_hd__nand2_1 _38999_ (.A(_16631_),
    .B(_15758_),
    .Y(_16632_));
 sky130_fd_sc_hd__and3_1 _39000_ (.A(_16626_),
    .B(_16629_),
    .C(_16627_),
    .X(_16633_));
 sky130_fd_sc_hd__o21ai_2 _39001_ (.A1(_16630_),
    .A2(_16633_),
    .B1(_15755_),
    .Y(_16634_));
 sky130_fd_sc_hd__nand2_1 _39002_ (.A(_16427_),
    .B(_16424_),
    .Y(_16635_));
 sky130_fd_sc_hd__o211ai_4 _39003_ (.A1(_16630_),
    .A2(_16632_),
    .B1(_16634_),
    .C1(_16635_),
    .Y(_16636_));
 sky130_fd_sc_hd__o21ai_2 _39004_ (.A1(_16630_),
    .A2(_16633_),
    .B1(_15758_),
    .Y(_16637_));
 sky130_fd_sc_hd__a21boi_2 _39005_ (.A1(_16423_),
    .A2(_16425_),
    .B1_N(_16424_),
    .Y(_16638_));
 sky130_fd_sc_hd__a21o_1 _39006_ (.A1(_16626_),
    .A2(_16627_),
    .B1(_16629_),
    .X(_16639_));
 sky130_fd_sc_hd__nand3_2 _39007_ (.A(_16639_),
    .B(_15755_),
    .C(_16631_),
    .Y(_16640_));
 sky130_fd_sc_hd__nand3_4 _39008_ (.A(_16637_),
    .B(_16638_),
    .C(_16640_),
    .Y(_16641_));
 sky130_vsdinv _39009_ (.A(_16456_),
    .Y(_16642_));
 sky130_fd_sc_hd__a21oi_2 _39010_ (.A1(_15758_),
    .A2(_16452_),
    .B1(_16642_),
    .Y(_16643_));
 sky130_vsdinv _39011_ (.A(_16643_),
    .Y(_16644_));
 sky130_fd_sc_hd__a21oi_4 _39012_ (.A1(_16636_),
    .A2(_16641_),
    .B1(_16644_),
    .Y(_16645_));
 sky130_fd_sc_hd__nand3_4 _39013_ (.A(_16636_),
    .B(_16641_),
    .C(_16644_),
    .Y(_16646_));
 sky130_vsdinv _39014_ (.A(_16646_),
    .Y(_16647_));
 sky130_fd_sc_hd__o2bb2ai_4 _39015_ (.A1_N(_16618_),
    .A2_N(_16622_),
    .B1(_16645_),
    .B2(_16647_),
    .Y(_16648_));
 sky130_fd_sc_hd__nor2_2 _39016_ (.A(_16645_),
    .B(_16647_),
    .Y(_16649_));
 sky130_fd_sc_hd__nand3_4 _39017_ (.A(_16649_),
    .B(_16618_),
    .C(_16622_),
    .Y(_16650_));
 sky130_fd_sc_hd__a21oi_2 _39018_ (.A1(_16429_),
    .A2(_16436_),
    .B1(_16430_),
    .Y(_16651_));
 sky130_fd_sc_hd__o21ai_4 _39019_ (.A1(_16472_),
    .A2(_16651_),
    .B1(_16437_),
    .Y(_16652_));
 sky130_fd_sc_hd__a21oi_4 _39020_ (.A1(_16648_),
    .A2(_16650_),
    .B1(_16652_),
    .Y(_16653_));
 sky130_fd_sc_hd__and3_1 _39021_ (.A(_16429_),
    .B(_16430_),
    .C(_16436_),
    .X(_16654_));
 sky130_fd_sc_hd__a31oi_1 _39022_ (.A1(_16439_),
    .A2(_16438_),
    .A3(_16440_),
    .B1(_16472_),
    .Y(_16655_));
 sky130_fd_sc_hd__o211a_2 _39023_ (.A1(_16654_),
    .A2(_16655_),
    .B1(_16650_),
    .C1(_16648_),
    .X(_16656_));
 sky130_fd_sc_hd__a21o_1 _39024_ (.A1(_16469_),
    .A2(_16464_),
    .B1(_16478_),
    .X(_16657_));
 sky130_fd_sc_hd__nand3_4 _39025_ (.A(_16478_),
    .B(_16469_),
    .C(_16464_),
    .Y(_16658_));
 sky130_fd_sc_hd__a21oi_4 _39026_ (.A1(_16657_),
    .A2(_16658_),
    .B1(_16484_),
    .Y(_16659_));
 sky130_fd_sc_hd__nand3_1 _39027_ (.A(_16657_),
    .B(_16482_),
    .C(_16658_),
    .Y(_16660_));
 sky130_vsdinv _39028_ (.A(_16660_),
    .Y(_16661_));
 sky130_fd_sc_hd__nor2_4 _39029_ (.A(_16659_),
    .B(_16661_),
    .Y(_16662_));
 sky130_fd_sc_hd__o21ai_4 _39030_ (.A1(_16653_),
    .A2(_16656_),
    .B1(_16662_),
    .Y(_16663_));
 sky130_fd_sc_hd__nand2_1 _39031_ (.A(_16491_),
    .B(_16490_),
    .Y(_16664_));
 sky130_fd_sc_hd__nand2_2 _39032_ (.A(_16664_),
    .B(_16489_),
    .Y(_16665_));
 sky130_fd_sc_hd__a21o_1 _39033_ (.A1(_16648_),
    .A2(_16650_),
    .B1(_16652_),
    .X(_16666_));
 sky130_fd_sc_hd__nand3_4 _39034_ (.A(_16652_),
    .B(_16650_),
    .C(_16648_),
    .Y(_16667_));
 sky130_fd_sc_hd__or2b_2 _39035_ (.A(_16659_),
    .B_N(_16660_),
    .X(_16668_));
 sky130_fd_sc_hd__nand3_4 _39036_ (.A(_16666_),
    .B(_16667_),
    .C(_16668_),
    .Y(_16669_));
 sky130_fd_sc_hd__nand3_4 _39037_ (.A(_16663_),
    .B(_16665_),
    .C(_16669_),
    .Y(_16670_));
 sky130_fd_sc_hd__o22ai_4 _39038_ (.A1(_16661_),
    .A2(_16659_),
    .B1(_16653_),
    .B2(_16656_),
    .Y(_16671_));
 sky130_fd_sc_hd__o21ai_2 _39039_ (.A1(_16490_),
    .A2(_16474_),
    .B1(_16491_),
    .Y(_16672_));
 sky130_fd_sc_hd__nand3_2 _39040_ (.A(_16666_),
    .B(_16667_),
    .C(_16662_),
    .Y(_16673_));
 sky130_fd_sc_hd__nand3_4 _39041_ (.A(_16671_),
    .B(_16672_),
    .C(_16673_),
    .Y(_16674_));
 sky130_fd_sc_hd__buf_6 _39042_ (.A(_14903_),
    .X(_16675_));
 sky130_fd_sc_hd__nand2_2 _39043_ (.A(_16485_),
    .B(_16477_),
    .Y(_16676_));
 sky130_fd_sc_hd__nor2_2 _39044_ (.A(_16675_),
    .B(_16676_),
    .Y(_16677_));
 sky130_vsdinv _39045_ (.A(_16676_),
    .Y(_16678_));
 sky130_fd_sc_hd__nor2_1 _39046_ (.A(_16313_),
    .B(_16678_),
    .Y(_16679_));
 sky130_fd_sc_hd__nor2_2 _39047_ (.A(_16677_),
    .B(_16679_),
    .Y(_16680_));
 sky130_fd_sc_hd__nand3_2 _39048_ (.A(_16670_),
    .B(_16674_),
    .C(_16680_),
    .Y(_16681_));
 sky130_fd_sc_hd__buf_2 _39049_ (.A(_16679_),
    .X(_16682_));
 sky130_fd_sc_hd__o2bb2ai_2 _39050_ (.A1_N(_16674_),
    .A2_N(_16670_),
    .B1(_16682_),
    .B2(_16677_),
    .Y(_16683_));
 sky130_fd_sc_hd__o211ai_4 _39051_ (.A1(_16532_),
    .A2(_16533_),
    .B1(_16681_),
    .C1(_16683_),
    .Y(_16684_));
 sky130_fd_sc_hd__a21boi_2 _39052_ (.A1(_16493_),
    .A2(_16502_),
    .B1_N(_16497_),
    .Y(_16685_));
 sky130_fd_sc_hd__nor2_4 _39053_ (.A(_16675_),
    .B(_16678_),
    .Y(_16686_));
 sky130_fd_sc_hd__nor2_4 _39054_ (.A(_14330_),
    .B(_16676_),
    .Y(_16687_));
 sky130_fd_sc_hd__o2bb2ai_2 _39055_ (.A1_N(_16674_),
    .A2_N(_16670_),
    .B1(_16686_),
    .B2(_16687_),
    .Y(_16688_));
 sky130_fd_sc_hd__nor2_4 _39056_ (.A(_16687_),
    .B(_16686_),
    .Y(_16689_));
 sky130_fd_sc_hd__nand3_2 _39057_ (.A(_16670_),
    .B(_16674_),
    .C(_16689_),
    .Y(_16690_));
 sky130_fd_sc_hd__nand3_4 _39058_ (.A(_16685_),
    .B(_16688_),
    .C(_16690_),
    .Y(_16691_));
 sky130_fd_sc_hd__nor2_8 _39059_ (.A(net410),
    .B(_16500_),
    .Y(_16692_));
 sky130_fd_sc_hd__nand3_4 _39060_ (.A(_16684_),
    .B(_16691_),
    .C(_16692_),
    .Y(_16693_));
 sky130_fd_sc_hd__nand2_1 _39061_ (.A(_16512_),
    .B(_16316_),
    .Y(_16694_));
 sky130_fd_sc_hd__a21oi_4 _39062_ (.A1(_16684_),
    .A2(_16691_),
    .B1(_16692_),
    .Y(_16695_));
 sky130_fd_sc_hd__a21oi_2 _39063_ (.A1(_16507_),
    .A2(_16694_),
    .B1(_16695_),
    .Y(_16696_));
 sky130_fd_sc_hd__nand2_2 _39064_ (.A(_16684_),
    .B(_16691_),
    .Y(_16697_));
 sky130_vsdinv _39065_ (.A(_16692_),
    .Y(_16698_));
 sky130_fd_sc_hd__nand2_1 _39066_ (.A(_16697_),
    .B(_16698_),
    .Y(_16699_));
 sky130_fd_sc_hd__nand2_1 _39067_ (.A(_16694_),
    .B(_16507_),
    .Y(_16700_));
 sky130_fd_sc_hd__a21oi_4 _39068_ (.A1(_16699_),
    .A2(_16693_),
    .B1(_16700_),
    .Y(_16701_));
 sky130_fd_sc_hd__a21oi_4 _39069_ (.A1(_16693_),
    .A2(_16696_),
    .B1(_16701_),
    .Y(_16702_));
 sky130_vsdinv _39070_ (.A(_16524_),
    .Y(_16703_));
 sky130_fd_sc_hd__nand3_4 _39071_ (.A(_16516_),
    .B(_16518_),
    .C(_16513_),
    .Y(_16704_));
 sky130_fd_sc_hd__o21ai_4 _39072_ (.A1(_16703_),
    .A2(_16531_),
    .B1(_16704_),
    .Y(_16705_));
 sky130_fd_sc_hd__xor2_4 _39073_ (.A(_16702_),
    .B(_16705_),
    .X(_02670_));
 sky130_fd_sc_hd__a31oi_4 _39074_ (.A1(_16663_),
    .A2(_16665_),
    .A3(_16669_),
    .B1(_16689_),
    .Y(_16706_));
 sky130_vsdinv _39075_ (.A(_16674_),
    .Y(_16707_));
 sky130_fd_sc_hd__nand2_1 _39076_ (.A(_16627_),
    .B(_16623_),
    .Y(_16708_));
 sky130_fd_sc_hd__nand2_2 _39077_ (.A(_16257_),
    .B(_19642_),
    .Y(_16709_));
 sky130_fd_sc_hd__o21ai_1 _39078_ (.A1(_15729_),
    .A2(_16258_),
    .B1(_16709_),
    .Y(_16710_));
 sky130_vsdinv _39079_ (.A(_16413_),
    .Y(_16711_));
 sky130_fd_sc_hd__o21bai_2 _39080_ (.A1(_16599_),
    .A2(_16711_),
    .B1_N(_16597_),
    .Y(_16712_));
 sky130_fd_sc_hd__xnor2_1 _39081_ (.A(_16710_),
    .B(_16712_),
    .Y(_16713_));
 sky130_fd_sc_hd__nand2_2 _39082_ (.A(_16708_),
    .B(_16713_),
    .Y(_16714_));
 sky130_fd_sc_hd__nand3b_4 _39083_ (.A_N(_16713_),
    .B(_16627_),
    .C(_16623_),
    .Y(_16715_));
 sky130_fd_sc_hd__a21o_1 _39084_ (.A1(_16714_),
    .A2(_16715_),
    .B1(_15754_),
    .X(_16716_));
 sky130_fd_sc_hd__nand3_4 _39085_ (.A(_16714_),
    .B(_15754_),
    .C(_16715_),
    .Y(_16717_));
 sky130_fd_sc_hd__nand2_1 _39086_ (.A(_16716_),
    .B(_16717_),
    .Y(_16718_));
 sky130_vsdinv _39087_ (.A(_16608_),
    .Y(_16719_));
 sky130_fd_sc_hd__a21oi_2 _39088_ (.A1(_16602_),
    .A2(_16603_),
    .B1(_16605_),
    .Y(_16720_));
 sky130_fd_sc_hd__o21ai_4 _39089_ (.A1(_16719_),
    .A2(_16720_),
    .B1(_16607_),
    .Y(_16721_));
 sky130_fd_sc_hd__nand2_4 _39090_ (.A(_16718_),
    .B(_16721_),
    .Y(_16722_));
 sky130_fd_sc_hd__nand3b_4 _39091_ (.A_N(_16721_),
    .B(_16716_),
    .C(_16717_),
    .Y(_16723_));
 sky130_fd_sc_hd__nand2_1 _39092_ (.A(_16722_),
    .B(_16723_),
    .Y(_16724_));
 sky130_fd_sc_hd__a21oi_2 _39093_ (.A1(_16639_),
    .A2(_15758_),
    .B1(_16633_),
    .Y(_16725_));
 sky130_fd_sc_hd__nand2_1 _39094_ (.A(_16724_),
    .B(_16725_),
    .Y(_16726_));
 sky130_vsdinv _39095_ (.A(_16726_),
    .Y(_16727_));
 sky130_vsdinv _39096_ (.A(_16725_),
    .Y(_16728_));
 sky130_fd_sc_hd__nand3_4 _39097_ (.A(_16722_),
    .B(_16723_),
    .C(_16728_),
    .Y(_16729_));
 sky130_vsdinv _39098_ (.A(_16729_),
    .Y(_16730_));
 sky130_fd_sc_hd__a21oi_4 _39099_ (.A1(_16558_),
    .A2(_16561_),
    .B1(_16559_),
    .Y(_16731_));
 sky130_fd_sc_hd__a21o_1 _39100_ (.A1(_16577_),
    .A2(_16562_),
    .B1(_16731_),
    .X(_16732_));
 sky130_fd_sc_hd__nor2_4 _39101_ (.A(_15814_),
    .B(_12078_),
    .Y(_16733_));
 sky130_fd_sc_hd__and4_2 _39102_ (.A(_10654_),
    .B(_13107_),
    .C(_19577_),
    .D(_10738_),
    .X(_16734_));
 sky130_fd_sc_hd__o22a_2 _39103_ (.A1(_11724_),
    .A2(_13745_),
    .B1(_15939_),
    .B2(_09765_),
    .X(_16735_));
 sky130_fd_sc_hd__nor2_2 _39104_ (.A(_16734_),
    .B(_16735_),
    .Y(_16736_));
 sky130_fd_sc_hd__nor2_2 _39105_ (.A(_16733_),
    .B(_16736_),
    .Y(_16737_));
 sky130_vsdinv _39106_ (.A(_16737_),
    .Y(_16738_));
 sky130_fd_sc_hd__nor2_1 _39107_ (.A(_16534_),
    .B(_16535_),
    .Y(_16739_));
 sky130_fd_sc_hd__nor2_2 _39108_ (.A(_16536_),
    .B(_16739_),
    .Y(_16740_));
 sky130_fd_sc_hd__nand2_2 _39109_ (.A(_16736_),
    .B(_16733_),
    .Y(_16741_));
 sky130_fd_sc_hd__nand3_4 _39110_ (.A(_16738_),
    .B(_16740_),
    .C(_16741_),
    .Y(_16742_));
 sky130_vsdinv _39111_ (.A(_16741_),
    .Y(_16743_));
 sky130_fd_sc_hd__o21bai_4 _39112_ (.A1(_16737_),
    .A2(_16743_),
    .B1_N(_16740_),
    .Y(_16744_));
 sky130_fd_sc_hd__a22o_1 _39113_ (.A1(_19583_),
    .A2(_19859_),
    .B1(_19588_),
    .B2(_19855_),
    .X(_16745_));
 sky130_fd_sc_hd__o31a_1 _39114_ (.A1(_15928_),
    .A2(_09929_),
    .A3(_15802_),
    .B1(_16745_),
    .X(_16746_));
 sky130_fd_sc_hd__nor2_4 _39115_ (.A(net468),
    .B(_13855_),
    .Y(_16747_));
 sky130_fd_sc_hd__and2_4 _39116_ (.A(_16746_),
    .B(_16747_),
    .X(_16748_));
 sky130_fd_sc_hd__nor2_4 _39117_ (.A(_16747_),
    .B(_16746_),
    .Y(_16749_));
 sky130_fd_sc_hd__o2bb2ai_4 _39118_ (.A1_N(_16742_),
    .A2_N(_16744_),
    .B1(_16748_),
    .B2(_16749_),
    .Y(_16750_));
 sky130_fd_sc_hd__nor2_4 _39119_ (.A(_16749_),
    .B(_16748_),
    .Y(_16751_));
 sky130_fd_sc_hd__nand3_4 _39120_ (.A(_16744_),
    .B(_16742_),
    .C(_16751_),
    .Y(_16752_));
 sky130_fd_sc_hd__nand2_4 _39121_ (.A(_16552_),
    .B(_16560_),
    .Y(_16753_));
 sky130_fd_sc_hd__a21oi_4 _39122_ (.A1(_16750_),
    .A2(_16752_),
    .B1(_16753_),
    .Y(_16754_));
 sky130_fd_sc_hd__a31oi_1 _39123_ (.A1(_16538_),
    .A2(_16540_),
    .A3(_16537_),
    .B1(_16554_),
    .Y(_16755_));
 sky130_fd_sc_hd__o211a_2 _39124_ (.A1(_16541_),
    .A2(_16755_),
    .B1(_16752_),
    .C1(_16750_),
    .X(_16756_));
 sky130_fd_sc_hd__and2b_2 _39125_ (.A_N(_16563_),
    .B(_16567_),
    .X(_16757_));
 sky130_fd_sc_hd__nand2_2 _39126_ (.A(_19597_),
    .B(_11228_),
    .Y(_16758_));
 sky130_fd_sc_hd__nand2_2 _39127_ (.A(_19600_),
    .B(_09950_),
    .Y(_16759_));
 sky130_fd_sc_hd__nor2_1 _39128_ (.A(_16758_),
    .B(_16759_),
    .Y(_16760_));
 sky130_fd_sc_hd__and2_1 _39129_ (.A(_16758_),
    .B(_16759_),
    .X(_16761_));
 sky130_fd_sc_hd__or4_4 _39130_ (.A(_08580_),
    .B(_12902_),
    .C(_16760_),
    .D(_16761_),
    .X(_16762_));
 sky130_fd_sc_hd__a2bb2o_2 _39131_ (.A1_N(_16760_),
    .A2_N(_16761_),
    .B1(_19604_),
    .B2(_19841_),
    .X(_16763_));
 sky130_fd_sc_hd__o21bai_4 _39132_ (.A1(_16544_),
    .A2(_16542_),
    .B1_N(_16546_),
    .Y(_16764_));
 sky130_fd_sc_hd__a21oi_4 _39133_ (.A1(_16762_),
    .A2(_16763_),
    .B1(_16764_),
    .Y(_16765_));
 sky130_fd_sc_hd__nor2_2 _39134_ (.A(_16757_),
    .B(_16765_),
    .Y(_16766_));
 sky130_fd_sc_hd__nand3_4 _39135_ (.A(_16762_),
    .B(_16764_),
    .C(_16763_),
    .Y(_16767_));
 sky130_fd_sc_hd__nand2_1 _39136_ (.A(_16766_),
    .B(_16767_),
    .Y(_16768_));
 sky130_vsdinv _39137_ (.A(_16767_),
    .Y(_16769_));
 sky130_fd_sc_hd__o21ai_1 _39138_ (.A1(_16765_),
    .A2(_16769_),
    .B1(_16757_),
    .Y(_16770_));
 sky130_fd_sc_hd__nand2_1 _39139_ (.A(_16768_),
    .B(_16770_),
    .Y(_16771_));
 sky130_fd_sc_hd__clkbuf_4 _39140_ (.A(_16771_),
    .X(_16772_));
 sky130_fd_sc_hd__o21ai_2 _39141_ (.A1(_16754_),
    .A2(_16756_),
    .B1(_16772_),
    .Y(_16773_));
 sky130_fd_sc_hd__a21o_1 _39142_ (.A1(_16750_),
    .A2(_16752_),
    .B1(_16753_),
    .X(_16774_));
 sky130_fd_sc_hd__nand3_4 _39143_ (.A(_16753_),
    .B(_16750_),
    .C(_16752_),
    .Y(_16775_));
 sky130_fd_sc_hd__nand3b_4 _39144_ (.A_N(_16772_),
    .B(_16774_),
    .C(_16775_),
    .Y(_16776_));
 sky130_fd_sc_hd__nand3_4 _39145_ (.A(_16732_),
    .B(_16773_),
    .C(_16776_),
    .Y(_16777_));
 sky130_fd_sc_hd__o21bai_4 _39146_ (.A1(_16754_),
    .A2(_16756_),
    .B1_N(_16772_),
    .Y(_16778_));
 sky130_fd_sc_hd__a21oi_4 _39147_ (.A1(_16577_),
    .A2(_16562_),
    .B1(_16731_),
    .Y(_16779_));
 sky130_fd_sc_hd__nand3_4 _39148_ (.A(_16774_),
    .B(_16775_),
    .C(_16772_),
    .Y(_16780_));
 sky130_fd_sc_hd__nand3_4 _39149_ (.A(_16778_),
    .B(_16779_),
    .C(_16780_),
    .Y(_16781_));
 sky130_fd_sc_hd__nand2_4 _39150_ (.A(_12274_),
    .B(_07822_),
    .Y(_16782_));
 sky130_fd_sc_hd__or2b_4 _39151_ (.A(_16782_),
    .B_N(_07758_),
    .X(_16783_));
 sky130_fd_sc_hd__nand2_2 _39152_ (.A(_16598_),
    .B(_16782_),
    .Y(_16784_));
 sky130_fd_sc_hd__nand2_1 _39153_ (.A(_16783_),
    .B(_16784_),
    .Y(_16785_));
 sky130_fd_sc_hd__or2_1 _39154_ (.A(_16711_),
    .B(_16785_),
    .X(_16786_));
 sky130_fd_sc_hd__buf_2 _39155_ (.A(_16786_),
    .X(_16787_));
 sky130_fd_sc_hd__nand2_2 _39156_ (.A(_16785_),
    .B(_16711_),
    .Y(_16788_));
 sky130_fd_sc_hd__nand2_2 _39157_ (.A(_15769_),
    .B(_19835_),
    .Y(_16789_));
 sky130_fd_sc_hd__nand2_2 _39158_ (.A(_15768_),
    .B(_19830_),
    .Y(_16790_));
 sky130_fd_sc_hd__or2_4 _39159_ (.A(_16789_),
    .B(_16790_),
    .X(_16791_));
 sky130_fd_sc_hd__nand2_2 _39160_ (.A(_16789_),
    .B(_16790_),
    .Y(_16792_));
 sky130_fd_sc_hd__nand2_1 _39161_ (.A(_16791_),
    .B(_16792_),
    .Y(_16793_));
 sky130_fd_sc_hd__nand2_2 _39162_ (.A(_19618_),
    .B(_19826_),
    .Y(_16794_));
 sky130_fd_sc_hd__nand2_2 _39163_ (.A(_16793_),
    .B(_16794_),
    .Y(_16795_));
 sky130_fd_sc_hd__nand3b_4 _39164_ (.A_N(_16794_),
    .B(_16791_),
    .C(_16792_),
    .Y(_16796_));
 sky130_fd_sc_hd__o21bai_2 _39165_ (.A1(_16587_),
    .A2(_16591_),
    .B1_N(_16590_),
    .Y(_16797_));
 sky130_fd_sc_hd__a21o_1 _39166_ (.A1(_16795_),
    .A2(_16796_),
    .B1(_16797_),
    .X(_16798_));
 sky130_fd_sc_hd__nand3_4 _39167_ (.A(_16795_),
    .B(_16797_),
    .C(_16796_),
    .Y(_16799_));
 sky130_fd_sc_hd__a22o_1 _39168_ (.A1(_16787_),
    .A2(_16788_),
    .B1(_16798_),
    .B2(_16799_),
    .X(_16800_));
 sky130_fd_sc_hd__and2_1 _39169_ (.A(_16786_),
    .B(_16788_),
    .X(_16801_));
 sky130_fd_sc_hd__buf_6 _39170_ (.A(_16801_),
    .X(_16802_));
 sky130_fd_sc_hd__nand3_4 _39171_ (.A(_16802_),
    .B(_16798_),
    .C(_16799_),
    .Y(_16803_));
 sky130_vsdinv _39172_ (.A(_16571_),
    .Y(_16804_));
 sky130_fd_sc_hd__o21ai_2 _39173_ (.A1(_16804_),
    .A2(_16572_),
    .B1(_16574_),
    .Y(_16805_));
 sky130_fd_sc_hd__a21o_1 _39174_ (.A1(_16800_),
    .A2(_16803_),
    .B1(_16805_),
    .X(_16806_));
 sky130_fd_sc_hd__nand3_4 _39175_ (.A(_16805_),
    .B(_16800_),
    .C(_16803_),
    .Y(_16807_));
 sky130_fd_sc_hd__nand2_1 _39176_ (.A(_16806_),
    .B(_16807_),
    .Y(_16808_));
 sky130_fd_sc_hd__nand2_2 _39177_ (.A(_16603_),
    .B(_16596_),
    .Y(_16809_));
 sky130_vsdinv _39178_ (.A(_16809_),
    .Y(_16810_));
 sky130_fd_sc_hd__nand2_1 _39179_ (.A(_16808_),
    .B(_16810_),
    .Y(_16811_));
 sky130_fd_sc_hd__nand3_4 _39180_ (.A(_16806_),
    .B(_16809_),
    .C(_16807_),
    .Y(_16812_));
 sky130_fd_sc_hd__and2_1 _39181_ (.A(_16811_),
    .B(_16812_),
    .X(_16813_));
 sky130_fd_sc_hd__a21o_2 _39182_ (.A1(_16777_),
    .A2(_16781_),
    .B1(_16813_),
    .X(_16814_));
 sky130_fd_sc_hd__nand3_4 _39183_ (.A(_16813_),
    .B(_16777_),
    .C(_16781_),
    .Y(_16815_));
 sky130_fd_sc_hd__o21ai_4 _39184_ (.A1(_16611_),
    .A2(_16582_),
    .B1(_16615_),
    .Y(_16816_));
 sky130_fd_sc_hd__a21oi_4 _39185_ (.A1(_16814_),
    .A2(_16815_),
    .B1(_16816_),
    .Y(_16817_));
 sky130_fd_sc_hd__and3_1 _39186_ (.A(_16732_),
    .B(_16773_),
    .C(_16776_),
    .X(_16818_));
 sky130_fd_sc_hd__nand2_1 _39187_ (.A(_16813_),
    .B(_16781_),
    .Y(_16819_));
 sky130_fd_sc_hd__o211a_1 _39188_ (.A1(_16818_),
    .A2(_16819_),
    .B1(_16814_),
    .C1(_16816_),
    .X(_16820_));
 sky130_fd_sc_hd__o22ai_4 _39189_ (.A1(_16727_),
    .A2(_16730_),
    .B1(_16817_),
    .B2(_16820_),
    .Y(_16821_));
 sky130_fd_sc_hd__nand2_2 _39190_ (.A(_16726_),
    .B(_16729_),
    .Y(_16822_));
 sky130_fd_sc_hd__a21o_1 _39191_ (.A1(_16814_),
    .A2(_16815_),
    .B1(_16816_),
    .X(_16823_));
 sky130_fd_sc_hd__nand3_4 _39192_ (.A(_16816_),
    .B(_16814_),
    .C(_16815_),
    .Y(_16824_));
 sky130_fd_sc_hd__nand3b_4 _39193_ (.A_N(_16822_),
    .B(_16823_),
    .C(_16824_),
    .Y(_16825_));
 sky130_fd_sc_hd__nand2_1 _39194_ (.A(_16649_),
    .B(_16622_),
    .Y(_16826_));
 sky130_fd_sc_hd__nand2_4 _39195_ (.A(_16826_),
    .B(_16618_),
    .Y(_16827_));
 sky130_fd_sc_hd__a21oi_4 _39196_ (.A1(_16821_),
    .A2(_16825_),
    .B1(_16827_),
    .Y(_16828_));
 sky130_vsdinv _39197_ (.A(_16618_),
    .Y(_16829_));
 sky130_fd_sc_hd__nand2_1 _39198_ (.A(_16636_),
    .B(_16641_),
    .Y(_16830_));
 sky130_fd_sc_hd__nand2_1 _39199_ (.A(_16830_),
    .B(_16643_),
    .Y(_16831_));
 sky130_fd_sc_hd__nand2_1 _39200_ (.A(_16831_),
    .B(_16646_),
    .Y(_16832_));
 sky130_fd_sc_hd__a31oi_1 _39201_ (.A1(_16620_),
    .A2(_16619_),
    .A3(_16621_),
    .B1(_16832_),
    .Y(_16833_));
 sky130_fd_sc_hd__o211a_1 _39202_ (.A1(_16829_),
    .A2(_16833_),
    .B1(_16825_),
    .C1(_16821_),
    .X(_16834_));
 sky130_fd_sc_hd__buf_4 _39203_ (.A(_16147_),
    .X(_16835_));
 sky130_fd_sc_hd__nand2_4 _39204_ (.A(_16646_),
    .B(_16636_),
    .Y(_16836_));
 sky130_fd_sc_hd__nor2_8 _39205_ (.A(_16835_),
    .B(_16836_),
    .Y(_16837_));
 sky130_fd_sc_hd__nand2_2 _39206_ (.A(_16836_),
    .B(_16835_),
    .Y(_16838_));
 sky130_fd_sc_hd__nand2_2 _39207_ (.A(_16838_),
    .B(_16482_),
    .Y(_16839_));
 sky130_fd_sc_hd__and2_1 _39208_ (.A(_16836_),
    .B(_16147_),
    .X(_16840_));
 sky130_vsdinv _39209_ (.A(_16481_),
    .Y(_16841_));
 sky130_fd_sc_hd__o21ai_2 _39210_ (.A1(_16837_),
    .A2(_16840_),
    .B1(_16841_),
    .Y(_16842_));
 sky130_fd_sc_hd__o21a_1 _39211_ (.A1(_16837_),
    .A2(_16839_),
    .B1(_16842_),
    .X(_16843_));
 sky130_fd_sc_hd__o21ai_2 _39212_ (.A1(_16828_),
    .A2(_16834_),
    .B1(_16843_),
    .Y(_16844_));
 sky130_fd_sc_hd__a21oi_2 _39213_ (.A1(_16666_),
    .A2(_16662_),
    .B1(_16656_),
    .Y(_16845_));
 sky130_fd_sc_hd__a21o_1 _39214_ (.A1(_16821_),
    .A2(_16825_),
    .B1(_16827_),
    .X(_16846_));
 sky130_fd_sc_hd__nand3_4 _39215_ (.A(_16827_),
    .B(_16821_),
    .C(_16825_),
    .Y(_16847_));
 sky130_fd_sc_hd__o21ai_2 _39216_ (.A1(_16837_),
    .A2(_16839_),
    .B1(_16842_),
    .Y(_16848_));
 sky130_fd_sc_hd__nand3_2 _39217_ (.A(_16846_),
    .B(_16847_),
    .C(_16848_),
    .Y(_16849_));
 sky130_fd_sc_hd__nand3_4 _39218_ (.A(_16844_),
    .B(_16845_),
    .C(_16849_),
    .Y(_16850_));
 sky130_fd_sc_hd__nor2_4 _39219_ (.A(_16837_),
    .B(_16839_),
    .Y(_16851_));
 sky130_vsdinv _39220_ (.A(_16842_),
    .Y(_16852_));
 sky130_fd_sc_hd__o22ai_4 _39221_ (.A1(_16851_),
    .A2(_16852_),
    .B1(_16828_),
    .B2(_16834_),
    .Y(_16853_));
 sky130_fd_sc_hd__nand3_2 _39222_ (.A(_16846_),
    .B(_16847_),
    .C(_16843_),
    .Y(_16854_));
 sky130_fd_sc_hd__o21ai_2 _39223_ (.A1(_16668_),
    .A2(_16653_),
    .B1(_16667_),
    .Y(_16855_));
 sky130_fd_sc_hd__nand3_4 _39224_ (.A(_16853_),
    .B(_16854_),
    .C(_16855_),
    .Y(_16856_));
 sky130_fd_sc_hd__nand2_1 _39225_ (.A(_16658_),
    .B(_16484_),
    .Y(_16857_));
 sky130_fd_sc_hd__nand2_2 _39226_ (.A(_16857_),
    .B(_16657_),
    .Y(_16858_));
 sky130_fd_sc_hd__nor2_4 _39227_ (.A(_16317_),
    .B(_16858_),
    .Y(_16859_));
 sky130_fd_sc_hd__nand2_1 _39228_ (.A(_16858_),
    .B(_14903_),
    .Y(_16860_));
 sky130_vsdinv _39229_ (.A(_16860_),
    .Y(_16861_));
 sky130_fd_sc_hd__nor2_4 _39230_ (.A(_16859_),
    .B(_16861_),
    .Y(_16862_));
 sky130_fd_sc_hd__nand3_2 _39231_ (.A(_16850_),
    .B(_16856_),
    .C(_16862_),
    .Y(_16863_));
 sky130_fd_sc_hd__buf_2 _39232_ (.A(_16861_),
    .X(_16864_));
 sky130_fd_sc_hd__o2bb2ai_2 _39233_ (.A1_N(_16856_),
    .A2_N(_16850_),
    .B1(_16864_),
    .B2(_16859_),
    .Y(_16865_));
 sky130_fd_sc_hd__o211ai_4 _39234_ (.A1(_16706_),
    .A2(_16707_),
    .B1(_16863_),
    .C1(_16865_),
    .Y(_16866_));
 sky130_fd_sc_hd__nor2_1 _39235_ (.A(_14331_),
    .B(_16858_),
    .Y(_16867_));
 sky130_vsdinv _39236_ (.A(_16858_),
    .Y(_16868_));
 sky130_fd_sc_hd__nor2_1 _39237_ (.A(_16318_),
    .B(_16868_),
    .Y(_16869_));
 sky130_fd_sc_hd__o2bb2ai_2 _39238_ (.A1_N(_16856_),
    .A2_N(_16850_),
    .B1(_16867_),
    .B2(_16869_),
    .Y(_16870_));
 sky130_fd_sc_hd__a21boi_2 _39239_ (.A1(_16670_),
    .A2(_16680_),
    .B1_N(_16674_),
    .Y(_16871_));
 sky130_fd_sc_hd__nand3b_2 _39240_ (.A_N(_16862_),
    .B(_16850_),
    .C(_16856_),
    .Y(_16872_));
 sky130_fd_sc_hd__nand3_4 _39241_ (.A(_16870_),
    .B(_16871_),
    .C(_16872_),
    .Y(_16873_));
 sky130_fd_sc_hd__a21oi_2 _39242_ (.A1(_16866_),
    .A2(_16873_),
    .B1(_16682_),
    .Y(_16874_));
 sky130_fd_sc_hd__and3_1 _39243_ (.A(_16866_),
    .B(_16873_),
    .C(_16682_),
    .X(_16875_));
 sky130_fd_sc_hd__nand2_1 _39244_ (.A(_16691_),
    .B(_16692_),
    .Y(_16876_));
 sky130_fd_sc_hd__nand2_2 _39245_ (.A(_16876_),
    .B(_16684_),
    .Y(_16877_));
 sky130_fd_sc_hd__o21bai_4 _39246_ (.A1(_16874_),
    .A2(_16875_),
    .B1_N(_16877_),
    .Y(_16878_));
 sky130_fd_sc_hd__a21o_1 _39247_ (.A1(_16866_),
    .A2(_16873_),
    .B1(_16682_),
    .X(_16879_));
 sky130_fd_sc_hd__nand3_2 _39248_ (.A(_16866_),
    .B(_16873_),
    .C(_16682_),
    .Y(_16880_));
 sky130_fd_sc_hd__nand3_4 _39249_ (.A(_16879_),
    .B(_16877_),
    .C(_16880_),
    .Y(_16881_));
 sky130_fd_sc_hd__nand2_2 _39250_ (.A(_16878_),
    .B(_16881_),
    .Y(_16882_));
 sky130_fd_sc_hd__and3_2 _39251_ (.A(_16684_),
    .B(_16691_),
    .C(_16692_),
    .X(_16883_));
 sky130_fd_sc_hd__a21oi_2 _39252_ (.A1(_16508_),
    .A2(_16511_),
    .B1(_16509_),
    .Y(_16884_));
 sky130_fd_sc_hd__a31oi_4 _39253_ (.A1(_16508_),
    .A2(_16509_),
    .A3(_16511_),
    .B1(_16520_),
    .Y(_16885_));
 sky130_fd_sc_hd__o2bb2ai_4 _39254_ (.A1_N(_16698_),
    .A2_N(_16697_),
    .B1(_16884_),
    .B2(_16885_),
    .Y(_16886_));
 sky130_fd_sc_hd__o22ai_4 _39255_ (.A1(_16883_),
    .A2(_16886_),
    .B1(_16704_),
    .B2(_16701_),
    .Y(_16887_));
 sky130_fd_sc_hd__a31oi_4 _39256_ (.A1(_16530_),
    .A2(_16702_),
    .A3(_16525_),
    .B1(_16887_),
    .Y(_16888_));
 sky130_vsdinv _39257_ (.A(_16888_),
    .Y(_16889_));
 sky130_fd_sc_hd__o21bai_2 _39258_ (.A1(_16695_),
    .A2(_16883_),
    .B1_N(_16700_),
    .Y(_16890_));
 sky130_fd_sc_hd__o2111ai_4 _39259_ (.A1(_16883_),
    .A2(_16886_),
    .B1(_16524_),
    .C1(_16704_),
    .D1(_16890_),
    .Y(_16891_));
 sky130_fd_sc_hd__nor2_1 _39260_ (.A(_16891_),
    .B(_16527_),
    .Y(_16892_));
 sky130_fd_sc_hd__and2_2 _39261_ (.A(_16135_),
    .B(_16892_),
    .X(_16893_));
 sky130_fd_sc_hd__nor2_4 _39262_ (.A(_16889_),
    .B(_16893_),
    .Y(_16894_));
 sky130_fd_sc_hd__nor2_8 _39263_ (.A(_16882_),
    .B(_16894_),
    .Y(_16895_));
 sky130_fd_sc_hd__and2_2 _39264_ (.A(_16894_),
    .B(_16882_),
    .X(_16896_));
 sky130_fd_sc_hd__nor2_8 _39265_ (.A(_16895_),
    .B(_16896_),
    .Y(_02671_));
 sky130_fd_sc_hd__nand2_1 _39266_ (.A(_16812_),
    .B(_16807_),
    .Y(_16897_));
 sky130_fd_sc_hd__and2_1 _39267_ (.A(_16787_),
    .B(_16783_),
    .X(_16898_));
 sky130_fd_sc_hd__nor2_2 _39268_ (.A(_16258_),
    .B(_15729_),
    .Y(_16899_));
 sky130_fd_sc_hd__o21ai_1 _39269_ (.A1(_16899_),
    .A2(_16712_),
    .B1(_16709_),
    .Y(_16900_));
 sky130_fd_sc_hd__nand2_1 _39270_ (.A(_16898_),
    .B(_16900_),
    .Y(_16901_));
 sky130_fd_sc_hd__a21o_1 _39271_ (.A1(_16787_),
    .A2(_16783_),
    .B1(_16900_),
    .X(_16902_));
 sky130_fd_sc_hd__nand2_2 _39272_ (.A(_16901_),
    .B(_16902_),
    .Y(_16903_));
 sky130_fd_sc_hd__nor2_4 _39273_ (.A(_15748_),
    .B(_16903_),
    .Y(_16904_));
 sky130_fd_sc_hd__nand2_1 _39274_ (.A(_16903_),
    .B(_15748_),
    .Y(_16905_));
 sky130_vsdinv _39275_ (.A(_16905_),
    .Y(_16906_));
 sky130_fd_sc_hd__nor2_2 _39276_ (.A(_16904_),
    .B(_16906_),
    .Y(_16907_));
 sky130_fd_sc_hd__nand2_4 _39277_ (.A(_16897_),
    .B(_16907_),
    .Y(_16908_));
 sky130_fd_sc_hd__o211ai_4 _39278_ (.A1(_16904_),
    .A2(_16906_),
    .B1(_16807_),
    .C1(_16812_),
    .Y(_16909_));
 sky130_vsdinv _39279_ (.A(_16715_),
    .Y(_16910_));
 sky130_fd_sc_hd__o21ai_4 _39280_ (.A1(_16045_),
    .A2(_16910_),
    .B1(_16714_),
    .Y(_16911_));
 sky130_fd_sc_hd__a21oi_4 _39281_ (.A1(_16908_),
    .A2(_16909_),
    .B1(_16911_),
    .Y(_16912_));
 sky130_fd_sc_hd__nand3_4 _39282_ (.A(_16908_),
    .B(_16909_),
    .C(_16911_),
    .Y(_16913_));
 sky130_vsdinv _39283_ (.A(_16913_),
    .Y(_16914_));
 sky130_fd_sc_hd__nand2_2 _39284_ (.A(_16752_),
    .B(_16742_),
    .Y(_16915_));
 sky130_fd_sc_hd__and4_1 _39285_ (.A(_09765_),
    .B(_13107_),
    .C(_19577_),
    .D(_10981_),
    .X(_16916_));
 sky130_fd_sc_hd__o22a_2 _39286_ (.A1(_10745_),
    .A2(_18475_),
    .B1(_15939_),
    .B2(net439),
    .X(_16917_));
 sky130_fd_sc_hd__nor2_1 _39287_ (.A(_16916_),
    .B(_16917_),
    .Y(_16918_));
 sky130_fd_sc_hd__nor2_2 _39288_ (.A(_15823_),
    .B(_15802_),
    .Y(_16919_));
 sky130_fd_sc_hd__nand2_2 _39289_ (.A(_16918_),
    .B(_16919_),
    .Y(_16920_));
 sky130_fd_sc_hd__a21o_1 _39290_ (.A1(_19580_),
    .A2(_19860_),
    .B1(_16918_),
    .X(_16921_));
 sky130_fd_sc_hd__nor2_4 _39291_ (.A(_16733_),
    .B(_16734_),
    .Y(_16922_));
 sky130_fd_sc_hd__o2bb2ai_4 _39292_ (.A1_N(_16920_),
    .A2_N(_16921_),
    .B1(_16735_),
    .B2(_16922_),
    .Y(_16923_));
 sky130_fd_sc_hd__nor2_2 _39293_ (.A(_16735_),
    .B(_16922_),
    .Y(_16924_));
 sky130_fd_sc_hd__nand3_4 _39294_ (.A(_16921_),
    .B(_16920_),
    .C(_16924_),
    .Y(_16925_));
 sky130_fd_sc_hd__or3_4 _39295_ (.A(_15928_),
    .B(_11545_),
    .C(_10652_),
    .X(_16926_));
 sky130_fd_sc_hd__a22o_1 _39296_ (.A1(_19584_),
    .A2(_14501_),
    .B1(_19589_),
    .B2(_19852_),
    .X(_16927_));
 sky130_fd_sc_hd__nor2_1 _39297_ (.A(net468),
    .B(_13260_),
    .Y(_16928_));
 sky130_fd_sc_hd__a21o_1 _39298_ (.A1(_16926_),
    .A2(_16927_),
    .B1(_16928_),
    .X(_16929_));
 sky130_fd_sc_hd__nand3_2 _39299_ (.A(_16926_),
    .B(_16928_),
    .C(_16927_),
    .Y(_16930_));
 sky130_fd_sc_hd__and2_2 _39300_ (.A(_16929_),
    .B(_16930_),
    .X(_16931_));
 sky130_fd_sc_hd__a21o_1 _39301_ (.A1(_16923_),
    .A2(_16925_),
    .B1(_16931_),
    .X(_16932_));
 sky130_fd_sc_hd__nand3_4 _39302_ (.A(_16923_),
    .B(_16931_),
    .C(_16925_),
    .Y(_16933_));
 sky130_fd_sc_hd__nand3_4 _39303_ (.A(_16915_),
    .B(_16932_),
    .C(_16933_),
    .Y(_16934_));
 sky130_fd_sc_hd__a21oi_2 _39304_ (.A1(_16923_),
    .A2(_16925_),
    .B1(_16931_),
    .Y(_16935_));
 sky130_fd_sc_hd__and3_1 _39305_ (.A(_16923_),
    .B(_16931_),
    .C(_16925_),
    .X(_16936_));
 sky130_fd_sc_hd__a21boi_2 _39306_ (.A1(_16744_),
    .A2(_16751_),
    .B1_N(_16742_),
    .Y(_16937_));
 sky130_fd_sc_hd__o21ai_4 _39307_ (.A1(_16935_),
    .A2(_16936_),
    .B1(_16937_),
    .Y(_16938_));
 sky130_fd_sc_hd__and4_2 _39308_ (.A(_19598_),
    .B(_19601_),
    .C(_11574_),
    .D(_13248_),
    .X(_16939_));
 sky130_fd_sc_hd__clkbuf_2 _39309_ (.A(_15956_),
    .X(_16940_));
 sky130_fd_sc_hd__o22a_1 _39310_ (.A1(_16940_),
    .A2(_13900_),
    .B1(_16184_),
    .B2(_09805_),
    .X(_16941_));
 sky130_fd_sc_hd__nor2_4 _39311_ (.A(_16939_),
    .B(_16941_),
    .Y(_16942_));
 sky130_fd_sc_hd__a21o_1 _39312_ (.A1(_19605_),
    .A2(_19836_),
    .B1(_16942_),
    .X(_16943_));
 sky130_fd_sc_hd__nand3_4 _39313_ (.A(_16942_),
    .B(_19605_),
    .C(_19837_),
    .Y(_16944_));
 sky130_fd_sc_hd__nand2_1 _39314_ (.A(_16943_),
    .B(_16944_),
    .Y(_16945_));
 sky130_fd_sc_hd__clkbuf_2 _39315_ (.A(_15929_),
    .X(_16946_));
 sky130_fd_sc_hd__and3_1 _39316_ (.A(_16946_),
    .B(_19856_),
    .C(_19860_),
    .X(_16947_));
 sky130_fd_sc_hd__nor2_1 _39317_ (.A(_16947_),
    .B(_16748_),
    .Y(_16948_));
 sky130_fd_sc_hd__nand2_2 _39318_ (.A(_16945_),
    .B(_16948_),
    .Y(_16949_));
 sky130_fd_sc_hd__o211ai_4 _39319_ (.A1(_16947_),
    .A2(_16748_),
    .B1(_16944_),
    .C1(_16943_),
    .Y(_16950_));
 sky130_vsdinv _39320_ (.A(_16760_),
    .Y(_16951_));
 sky130_fd_sc_hd__nand2_2 _39321_ (.A(_16762_),
    .B(_16951_),
    .Y(_16952_));
 sky130_fd_sc_hd__nand3_2 _39322_ (.A(_16949_),
    .B(_16950_),
    .C(_16952_),
    .Y(_16953_));
 sky130_vsdinv _39323_ (.A(_16953_),
    .Y(_16954_));
 sky130_fd_sc_hd__nand2_1 _39324_ (.A(_16949_),
    .B(_16950_),
    .Y(_16955_));
 sky130_vsdinv _39325_ (.A(_16952_),
    .Y(_16956_));
 sky130_fd_sc_hd__nand2_1 _39326_ (.A(_16955_),
    .B(_16956_),
    .Y(_16957_));
 sky130_vsdinv _39327_ (.A(_16957_),
    .Y(_16958_));
 sky130_fd_sc_hd__o2bb2ai_4 _39328_ (.A1_N(_16934_),
    .A2_N(_16938_),
    .B1(_16954_),
    .B2(_16958_),
    .Y(_16959_));
 sky130_fd_sc_hd__nand2_2 _39329_ (.A(_16957_),
    .B(_16953_),
    .Y(_16960_));
 sky130_fd_sc_hd__nand3b_4 _39330_ (.A_N(_16960_),
    .B(_16938_),
    .C(_16934_),
    .Y(_16961_));
 sky130_fd_sc_hd__o21ai_4 _39331_ (.A1(_16772_),
    .A2(_16754_),
    .B1(_16775_),
    .Y(_16962_));
 sky130_fd_sc_hd__a21oi_4 _39332_ (.A1(_16959_),
    .A2(_16961_),
    .B1(_16962_),
    .Y(_16963_));
 sky130_fd_sc_hd__nor2_1 _39333_ (.A(_16772_),
    .B(_16754_),
    .Y(_16964_));
 sky130_fd_sc_hd__o211a_1 _39334_ (.A1(_16756_),
    .A2(_16964_),
    .B1(_16961_),
    .C1(_16959_),
    .X(_16965_));
 sky130_fd_sc_hd__nand2_1 _39335_ (.A(_15769_),
    .B(_11199_),
    .Y(_16966_));
 sky130_fd_sc_hd__nand2_2 _39336_ (.A(_12466_),
    .B(_11597_),
    .Y(_16967_));
 sky130_fd_sc_hd__or2_2 _39337_ (.A(_16966_),
    .B(_16967_),
    .X(_16968_));
 sky130_fd_sc_hd__nand2_1 _39338_ (.A(_16966_),
    .B(_16967_),
    .Y(_16969_));
 sky130_fd_sc_hd__nand2_4 _39339_ (.A(_11594_),
    .B(_19617_),
    .Y(_16970_));
 sky130_vsdinv _39340_ (.A(_16970_),
    .Y(_16971_));
 sky130_fd_sc_hd__a21o_1 _39341_ (.A1(_16968_),
    .A2(_16969_),
    .B1(_16971_),
    .X(_16972_));
 sky130_fd_sc_hd__nand3_2 _39342_ (.A(_16968_),
    .B(_16971_),
    .C(_16969_),
    .Y(_16973_));
 sky130_fd_sc_hd__nand2_2 _39343_ (.A(_16972_),
    .B(_16973_),
    .Y(_16974_));
 sky130_fd_sc_hd__a21o_1 _39344_ (.A1(_16791_),
    .A2(_16796_),
    .B1(_16974_),
    .X(_16975_));
 sky130_fd_sc_hd__nand3_4 _39345_ (.A(_16974_),
    .B(_16791_),
    .C(_16796_),
    .Y(_16976_));
 sky130_fd_sc_hd__nand2_4 _39346_ (.A(_16787_),
    .B(_16788_),
    .Y(_16977_));
 sky130_fd_sc_hd__a21o_1 _39347_ (.A1(_16975_),
    .A2(_16976_),
    .B1(_16977_),
    .X(_16978_));
 sky130_fd_sc_hd__nand3_4 _39348_ (.A(_16975_),
    .B(_16977_),
    .C(_16976_),
    .Y(_16979_));
 sky130_fd_sc_hd__o2bb2ai_4 _39349_ (.A1_N(_16978_),
    .A2_N(_16979_),
    .B1(_16769_),
    .B2(_16766_),
    .Y(_16980_));
 sky130_fd_sc_hd__o2111ai_4 _39350_ (.A1(_16757_),
    .A2(_16765_),
    .B1(_16767_),
    .C1(_16979_),
    .D1(_16978_),
    .Y(_16981_));
 sky130_fd_sc_hd__nand2_4 _39351_ (.A(_16803_),
    .B(_16799_),
    .Y(_16982_));
 sky130_fd_sc_hd__a21o_1 _39352_ (.A1(_16980_),
    .A2(_16981_),
    .B1(_16982_),
    .X(_16983_));
 sky130_fd_sc_hd__nand3_4 _39353_ (.A(_16980_),
    .B(_16982_),
    .C(_16981_),
    .Y(_16984_));
 sky130_fd_sc_hd__nand2_1 _39354_ (.A(_16983_),
    .B(_16984_),
    .Y(_16985_));
 sky130_fd_sc_hd__o21ai_2 _39355_ (.A1(_16963_),
    .A2(_16965_),
    .B1(_16985_),
    .Y(_16986_));
 sky130_fd_sc_hd__and2_1 _39356_ (.A(_16771_),
    .B(_16775_),
    .X(_16987_));
 sky130_fd_sc_hd__o2bb2ai_4 _39357_ (.A1_N(_16961_),
    .A2_N(_16959_),
    .B1(_16754_),
    .B2(_16987_),
    .Y(_16988_));
 sky130_fd_sc_hd__a21oi_4 _39358_ (.A1(_16980_),
    .A2(_16981_),
    .B1(_16982_),
    .Y(_16989_));
 sky130_fd_sc_hd__and3_2 _39359_ (.A(_16980_),
    .B(_16982_),
    .C(_16981_),
    .X(_16990_));
 sky130_fd_sc_hd__nor2_8 _39360_ (.A(_16989_),
    .B(_16990_),
    .Y(_16991_));
 sky130_fd_sc_hd__nand3_4 _39361_ (.A(_16959_),
    .B(_16962_),
    .C(_16961_),
    .Y(_16992_));
 sky130_fd_sc_hd__nand3_4 _39362_ (.A(_16988_),
    .B(_16991_),
    .C(_16992_),
    .Y(_16993_));
 sky130_fd_sc_hd__nand2_2 _39363_ (.A(_16819_),
    .B(_16777_),
    .Y(_16994_));
 sky130_fd_sc_hd__a21oi_4 _39364_ (.A1(_16986_),
    .A2(_16993_),
    .B1(_16994_),
    .Y(_16995_));
 sky130_fd_sc_hd__a21oi_4 _39365_ (.A1(_16988_),
    .A2(_16992_),
    .B1(_16991_),
    .Y(_16996_));
 sky130_fd_sc_hd__nand2_1 _39366_ (.A(_16811_),
    .B(_16812_),
    .Y(_16997_));
 sky130_fd_sc_hd__a31oi_4 _39367_ (.A1(_16779_),
    .A2(_16778_),
    .A3(_16780_),
    .B1(_16997_),
    .Y(_16998_));
 sky130_fd_sc_hd__o21ai_4 _39368_ (.A1(_16818_),
    .A2(_16998_),
    .B1(_16993_),
    .Y(_16999_));
 sky130_fd_sc_hd__nor2_2 _39369_ (.A(_16996_),
    .B(_16999_),
    .Y(_17000_));
 sky130_fd_sc_hd__o22ai_4 _39370_ (.A1(_16912_),
    .A2(_16914_),
    .B1(_16995_),
    .B2(_17000_),
    .Y(_17001_));
 sky130_fd_sc_hd__nor2_2 _39371_ (.A(_16912_),
    .B(_16914_),
    .Y(_17002_));
 sky130_fd_sc_hd__and3_1 _39372_ (.A(_16988_),
    .B(_16991_),
    .C(_16992_),
    .X(_17003_));
 sky130_fd_sc_hd__o21bai_2 _39373_ (.A1(_16996_),
    .A2(_17003_),
    .B1_N(_16994_),
    .Y(_17004_));
 sky130_fd_sc_hd__o211ai_4 _39374_ (.A1(_16996_),
    .A2(_16999_),
    .B1(_17002_),
    .C1(_17004_),
    .Y(_17005_));
 sky130_fd_sc_hd__o21ai_4 _39375_ (.A1(_16822_),
    .A2(_16817_),
    .B1(_16824_),
    .Y(_17006_));
 sky130_fd_sc_hd__a21oi_4 _39376_ (.A1(_17001_),
    .A2(_17005_),
    .B1(_17006_),
    .Y(_17007_));
 sky130_fd_sc_hd__nor2_1 _39377_ (.A(_16822_),
    .B(_16817_),
    .Y(_17008_));
 sky130_fd_sc_hd__o211a_1 _39378_ (.A1(_16820_),
    .A2(_17008_),
    .B1(_17005_),
    .C1(_17001_),
    .X(_17009_));
 sky130_fd_sc_hd__and2_1 _39379_ (.A(_16718_),
    .B(_16721_),
    .X(_17010_));
 sky130_fd_sc_hd__a211oi_4 _39380_ (.A1(_16723_),
    .A2(_16728_),
    .B1(_16835_),
    .C1(_17010_),
    .Y(_17011_));
 sky130_fd_sc_hd__clkbuf_4 _39381_ (.A(_16835_),
    .X(_17012_));
 sky130_fd_sc_hd__nand2_1 _39382_ (.A(_16729_),
    .B(_16722_),
    .Y(_17013_));
 sky130_fd_sc_hd__o2bb2ai_2 _39383_ (.A1_N(_17012_),
    .A2_N(_17013_),
    .B1(_16141_),
    .B2(_16144_),
    .Y(_17014_));
 sky130_fd_sc_hd__a21oi_4 _39384_ (.A1(_16729_),
    .A2(_16722_),
    .B1(_16478_),
    .Y(_17015_));
 sky130_fd_sc_hd__o22ai_4 _39385_ (.A1(_16145_),
    .A2(_16480_),
    .B1(_17011_),
    .B2(_17015_),
    .Y(_17016_));
 sky130_fd_sc_hd__o21a_2 _39386_ (.A1(_17011_),
    .A2(_17014_),
    .B1(_17016_),
    .X(_17017_));
 sky130_fd_sc_hd__o21ai_4 _39387_ (.A1(_17007_),
    .A2(_17009_),
    .B1(_17017_),
    .Y(_17018_));
 sky130_fd_sc_hd__nand2_1 _39388_ (.A(_16847_),
    .B(_16848_),
    .Y(_17019_));
 sky130_fd_sc_hd__nand2_4 _39389_ (.A(_17019_),
    .B(_16846_),
    .Y(_17020_));
 sky130_fd_sc_hd__a21o_2 _39390_ (.A1(_17001_),
    .A2(_17005_),
    .B1(_17006_),
    .X(_17021_));
 sky130_fd_sc_hd__nand3_4 _39391_ (.A(_17001_),
    .B(_17006_),
    .C(_17005_),
    .Y(_17022_));
 sky130_fd_sc_hd__o21ai_4 _39392_ (.A1(_17011_),
    .A2(_17014_),
    .B1(_17016_),
    .Y(_17023_));
 sky130_fd_sc_hd__nand3_4 _39393_ (.A(_17021_),
    .B(_17022_),
    .C(_17023_),
    .Y(_17024_));
 sky130_fd_sc_hd__nand3_4 _39394_ (.A(_17018_),
    .B(_17020_),
    .C(_17024_),
    .Y(_17025_));
 sky130_fd_sc_hd__o21ai_2 _39395_ (.A1(_17007_),
    .A2(_17009_),
    .B1(_17023_),
    .Y(_17026_));
 sky130_fd_sc_hd__o21ai_2 _39396_ (.A1(_16848_),
    .A2(_16828_),
    .B1(_16847_),
    .Y(_17027_));
 sky130_fd_sc_hd__nand3_4 _39397_ (.A(_17021_),
    .B(_17022_),
    .C(_17017_),
    .Y(_17028_));
 sky130_fd_sc_hd__nand3_4 _39398_ (.A(_17026_),
    .B(_17027_),
    .C(_17028_),
    .Y(_17029_));
 sky130_fd_sc_hd__nand2_1 _39399_ (.A(_17025_),
    .B(_17029_),
    .Y(_17030_));
 sky130_fd_sc_hd__or2_1 _39400_ (.A(_16841_),
    .B(_16837_),
    .X(_17031_));
 sky130_fd_sc_hd__nand2_4 _39401_ (.A(_17031_),
    .B(_16838_),
    .Y(_17032_));
 sky130_fd_sc_hd__nor2_4 _39402_ (.A(_16313_),
    .B(_17032_),
    .Y(_17033_));
 sky130_fd_sc_hd__nor2_2 _39403_ (.A(_16840_),
    .B(_16851_),
    .Y(_17034_));
 sky130_fd_sc_hd__nor2_4 _39404_ (.A(_16675_),
    .B(_17034_),
    .Y(_17035_));
 sky130_fd_sc_hd__nor2_4 _39405_ (.A(_17033_),
    .B(_17035_),
    .Y(_17036_));
 sky130_fd_sc_hd__nand2_2 _39406_ (.A(_17030_),
    .B(_17036_),
    .Y(_17037_));
 sky130_fd_sc_hd__nand2_1 _39407_ (.A(_16850_),
    .B(_16862_),
    .Y(_17038_));
 sky130_fd_sc_hd__nand2_2 _39408_ (.A(_17038_),
    .B(_16856_),
    .Y(_17039_));
 sky130_fd_sc_hd__nor2_4 _39409_ (.A(_16675_),
    .B(_17032_),
    .Y(_17040_));
 sky130_fd_sc_hd__nand2_2 _39410_ (.A(_17032_),
    .B(_16317_),
    .Y(_17041_));
 sky130_vsdinv _39411_ (.A(_17041_),
    .Y(_17042_));
 sky130_fd_sc_hd__nor2_8 _39412_ (.A(_17040_),
    .B(_17042_),
    .Y(_17043_));
 sky130_fd_sc_hd__nand3_4 _39413_ (.A(_17029_),
    .B(_17025_),
    .C(_17043_),
    .Y(_17044_));
 sky130_fd_sc_hd__nand3_4 _39414_ (.A(_17037_),
    .B(_17039_),
    .C(_17044_),
    .Y(_17045_));
 sky130_fd_sc_hd__o2bb2ai_2 _39415_ (.A1_N(_17025_),
    .A2_N(_17029_),
    .B1(_17033_),
    .B2(_17035_),
    .Y(_17046_));
 sky130_fd_sc_hd__a21boi_2 _39416_ (.A1(_16850_),
    .A2(_16862_),
    .B1_N(_16856_),
    .Y(_17047_));
 sky130_fd_sc_hd__nand3_2 _39417_ (.A(_17029_),
    .B(_17025_),
    .C(_17036_),
    .Y(_17048_));
 sky130_fd_sc_hd__nand3_4 _39418_ (.A(_17046_),
    .B(_17047_),
    .C(_17048_),
    .Y(_17049_));
 sky130_fd_sc_hd__a21oi_4 _39419_ (.A1(_17045_),
    .A2(_17049_),
    .B1(_16864_),
    .Y(_17050_));
 sky130_fd_sc_hd__and3_1 _39420_ (.A(_17045_),
    .B(_17049_),
    .C(_16864_),
    .X(_17051_));
 sky130_fd_sc_hd__nand2_1 _39421_ (.A(_16873_),
    .B(_16682_),
    .Y(_17052_));
 sky130_fd_sc_hd__nand2_2 _39422_ (.A(_17052_),
    .B(_16866_),
    .Y(_17053_));
 sky130_fd_sc_hd__o21bai_4 _39423_ (.A1(_17050_),
    .A2(_17051_),
    .B1_N(_17053_),
    .Y(_17054_));
 sky130_fd_sc_hd__a21o_1 _39424_ (.A1(_17045_),
    .A2(_17049_),
    .B1(_16864_),
    .X(_17055_));
 sky130_fd_sc_hd__nand3_2 _39425_ (.A(_17045_),
    .B(_17049_),
    .C(_16864_),
    .Y(_17056_));
 sky130_fd_sc_hd__nand3_1 _39426_ (.A(_17055_),
    .B(_17053_),
    .C(_17056_),
    .Y(_17057_));
 sky130_fd_sc_hd__and2_1 _39427_ (.A(_17054_),
    .B(_17057_),
    .X(_17058_));
 sky130_fd_sc_hd__nand3b_2 _39428_ (.A_N(_16895_),
    .B(_16881_),
    .C(_17058_),
    .Y(_17059_));
 sky130_vsdinv _39429_ (.A(_16881_),
    .Y(_17060_));
 sky130_fd_sc_hd__o21bai_2 _39430_ (.A1(_17060_),
    .A2(_16895_),
    .B1_N(_17058_),
    .Y(_17061_));
 sky130_fd_sc_hd__nand2_4 _39431_ (.A(_17059_),
    .B(_17061_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand2_2 _39432_ (.A(_17053_),
    .B(_17056_),
    .Y(_17062_));
 sky130_fd_sc_hd__o2111a_1 _39433_ (.A1(_17050_),
    .A2(_17062_),
    .B1(_16881_),
    .C1(_16878_),
    .D1(_17054_),
    .X(_17063_));
 sky130_fd_sc_hd__o21ai_1 _39434_ (.A1(_16889_),
    .A2(_16893_),
    .B1(_17063_),
    .Y(_17064_));
 sky130_fd_sc_hd__nand2_1 _39435_ (.A(_17057_),
    .B(_16881_),
    .Y(_17065_));
 sky130_fd_sc_hd__nand2_1 _39436_ (.A(_17065_),
    .B(_17054_),
    .Y(_17066_));
 sky130_fd_sc_hd__a21oi_4 _39437_ (.A1(_17018_),
    .A2(_17024_),
    .B1(_17020_),
    .Y(_17067_));
 sky130_fd_sc_hd__a31oi_4 _39438_ (.A1(_17018_),
    .A2(_17020_),
    .A3(_17024_),
    .B1(_17036_),
    .Y(_17068_));
 sky130_fd_sc_hd__a21oi_2 _39439_ (.A1(_16988_),
    .A2(_16991_),
    .B1(_16965_),
    .Y(_17069_));
 sky130_fd_sc_hd__nand2_2 _39440_ (.A(_16933_),
    .B(_16925_),
    .Y(_17070_));
 sky130_fd_sc_hd__nor2_8 _39441_ (.A(_15823_),
    .B(_09929_),
    .Y(_17071_));
 sky130_fd_sc_hd__and4_4 _39442_ (.A(net439),
    .B(_15937_),
    .C(_19577_),
    .D(_13413_),
    .X(_17072_));
 sky130_fd_sc_hd__o22a_4 _39443_ (.A1(_19864_),
    .A2(_18475_),
    .B1(_15939_),
    .B2(_15802_),
    .X(_17073_));
 sky130_fd_sc_hd__nor3_4 _39444_ (.A(_17071_),
    .B(_17072_),
    .C(_17073_),
    .Y(_17074_));
 sky130_fd_sc_hd__o21a_1 _39445_ (.A1(_17072_),
    .A2(_17073_),
    .B1(_17071_),
    .X(_17075_));
 sky130_fd_sc_hd__nor2_2 _39446_ (.A(_16919_),
    .B(_16916_),
    .Y(_17076_));
 sky130_fd_sc_hd__nor2_4 _39447_ (.A(_16917_),
    .B(_17076_),
    .Y(_17077_));
 sky130_fd_sc_hd__o21a_2 _39448_ (.A1(_17074_),
    .A2(_17075_),
    .B1(_17077_),
    .X(_17078_));
 sky130_fd_sc_hd__nor3_4 _39449_ (.A(_17074_),
    .B(_17075_),
    .C(_17077_),
    .Y(_17079_));
 sky130_fd_sc_hd__nand2_1 _39450_ (.A(_15806_),
    .B(_19845_),
    .Y(_17080_));
 sky130_vsdinv _39451_ (.A(_17080_),
    .Y(_17081_));
 sky130_fd_sc_hd__o22a_1 _39452_ (.A1(_16159_),
    .A2(_13855_),
    .B1(_15932_),
    .B2(_13260_),
    .X(_17082_));
 sky130_fd_sc_hd__and3_1 _39453_ (.A(_15929_),
    .B(_15316_),
    .C(_19852_),
    .X(_17083_));
 sky130_fd_sc_hd__nor2_4 _39454_ (.A(_17082_),
    .B(_17083_),
    .Y(_17084_));
 sky130_fd_sc_hd__or2_1 _39455_ (.A(_17081_),
    .B(_17084_),
    .X(_17085_));
 sky130_fd_sc_hd__nand2_1 _39456_ (.A(_17084_),
    .B(_17081_),
    .Y(_17086_));
 sky130_fd_sc_hd__nand2_2 _39457_ (.A(_17085_),
    .B(_17086_),
    .Y(_17087_));
 sky130_fd_sc_hd__o21ai_2 _39458_ (.A1(_17078_),
    .A2(_17079_),
    .B1(_17087_),
    .Y(_17088_));
 sky130_fd_sc_hd__nor2_1 _39459_ (.A(_17081_),
    .B(_17084_),
    .Y(_17089_));
 sky130_fd_sc_hd__and2b_1 _39460_ (.A_N(_17089_),
    .B(_17086_),
    .X(_17090_));
 sky130_vsdinv _39461_ (.A(_17079_),
    .Y(_17091_));
 sky130_vsdinv _39462_ (.A(_17078_),
    .Y(_17092_));
 sky130_fd_sc_hd__nand3_2 _39463_ (.A(_17090_),
    .B(_17091_),
    .C(_17092_),
    .Y(_17093_));
 sky130_fd_sc_hd__nand3_4 _39464_ (.A(_17070_),
    .B(_17088_),
    .C(_17093_),
    .Y(_17094_));
 sky130_fd_sc_hd__a21boi_2 _39465_ (.A1(_16923_),
    .A2(_16931_),
    .B1_N(_16925_),
    .Y(_17095_));
 sky130_fd_sc_hd__nand3_4 _39466_ (.A(_17091_),
    .B(_17087_),
    .C(_17092_),
    .Y(_17096_));
 sky130_fd_sc_hd__o21ai_2 _39467_ (.A1(_17078_),
    .A2(_17079_),
    .B1(_17090_),
    .Y(_17097_));
 sky130_fd_sc_hd__nand3_4 _39468_ (.A(_17095_),
    .B(_17096_),
    .C(_17097_),
    .Y(_17098_));
 sky130_fd_sc_hd__nor2_2 _39469_ (.A(_08580_),
    .B(_13309_),
    .Y(_17099_));
 sky130_fd_sc_hd__nand2_1 _39470_ (.A(_14087_),
    .B(_10601_),
    .Y(_17100_));
 sky130_fd_sc_hd__nand2_1 _39471_ (.A(_14084_),
    .B(_12639_),
    .Y(_17101_));
 sky130_fd_sc_hd__nor2_2 _39472_ (.A(_17100_),
    .B(_17101_),
    .Y(_17102_));
 sky130_fd_sc_hd__and2_1 _39473_ (.A(_17100_),
    .B(_17101_),
    .X(_17103_));
 sky130_fd_sc_hd__nor2_2 _39474_ (.A(_17102_),
    .B(_17103_),
    .Y(_17104_));
 sky130_fd_sc_hd__or2_2 _39475_ (.A(_17099_),
    .B(_17104_),
    .X(_17105_));
 sky130_fd_sc_hd__nand2_2 _39476_ (.A(_17104_),
    .B(_17099_),
    .Y(_17106_));
 sky130_fd_sc_hd__nand2_2 _39477_ (.A(_16930_),
    .B(_16926_),
    .Y(_17107_));
 sky130_fd_sc_hd__a21o_1 _39478_ (.A1(_17105_),
    .A2(_17106_),
    .B1(_17107_),
    .X(_17108_));
 sky130_fd_sc_hd__nand3_4 _39479_ (.A(_17107_),
    .B(_17105_),
    .C(_17106_),
    .Y(_17109_));
 sky130_fd_sc_hd__and3_1 _39480_ (.A(_16942_),
    .B(_19605_),
    .C(_19837_),
    .X(_17110_));
 sky130_fd_sc_hd__nor2_4 _39481_ (.A(_16939_),
    .B(_17110_),
    .Y(_17111_));
 sky130_fd_sc_hd__a21o_1 _39482_ (.A1(_17108_),
    .A2(_17109_),
    .B1(_17111_),
    .X(_17112_));
 sky130_fd_sc_hd__nand3_2 _39483_ (.A(_17108_),
    .B(_17111_),
    .C(_17109_),
    .Y(_17113_));
 sky130_fd_sc_hd__nand2_4 _39484_ (.A(_17112_),
    .B(_17113_),
    .Y(_17114_));
 sky130_fd_sc_hd__a21o_2 _39485_ (.A1(_17094_),
    .A2(_17098_),
    .B1(_17114_),
    .X(_17115_));
 sky130_fd_sc_hd__nand3_4 _39486_ (.A(_17094_),
    .B(_17114_),
    .C(_17098_),
    .Y(_17116_));
 sky130_fd_sc_hd__a21oi_2 _39487_ (.A1(_16932_),
    .A2(_16933_),
    .B1(_16915_),
    .Y(_17117_));
 sky130_fd_sc_hd__o21ai_4 _39488_ (.A1(_16960_),
    .A2(_17117_),
    .B1(_16934_),
    .Y(_17118_));
 sky130_fd_sc_hd__a21oi_4 _39489_ (.A1(_17115_),
    .A2(_17116_),
    .B1(_17118_),
    .Y(_17119_));
 sky130_vsdinv _39490_ (.A(_17094_),
    .Y(_17120_));
 sky130_fd_sc_hd__nand2_1 _39491_ (.A(_17114_),
    .B(_17098_),
    .Y(_17121_));
 sky130_fd_sc_hd__o211a_1 _39492_ (.A1(_17120_),
    .A2(_17121_),
    .B1(_17118_),
    .C1(_17115_),
    .X(_17122_));
 sky130_vsdinv _39493_ (.A(_16950_),
    .Y(_17123_));
 sky130_fd_sc_hd__a21o_1 _39494_ (.A1(_16952_),
    .A2(_16949_),
    .B1(_17123_),
    .X(_17124_));
 sky130_fd_sc_hd__nand2_2 _39495_ (.A(_19609_),
    .B(_19827_),
    .Y(_17125_));
 sky130_fd_sc_hd__nand2_4 _39496_ (.A(_11594_),
    .B(_15768_),
    .Y(_17126_));
 sky130_fd_sc_hd__xor2_4 _39497_ (.A(_16970_),
    .B(_17126_),
    .X(_17127_));
 sky130_fd_sc_hd__or2_1 _39498_ (.A(_17125_),
    .B(_17127_),
    .X(_17128_));
 sky130_fd_sc_hd__nand2_1 _39499_ (.A(_17127_),
    .B(_17125_),
    .Y(_17129_));
 sky130_fd_sc_hd__nand2_1 _39500_ (.A(_16973_),
    .B(_16968_),
    .Y(_17130_));
 sky130_vsdinv _39501_ (.A(_17130_),
    .Y(_17131_));
 sky130_fd_sc_hd__a21o_1 _39502_ (.A1(_17128_),
    .A2(_17129_),
    .B1(_17131_),
    .X(_17132_));
 sky130_fd_sc_hd__xor2_1 _39503_ (.A(_17125_),
    .B(_17127_),
    .X(_17133_));
 sky130_fd_sc_hd__nand2_1 _39504_ (.A(_17133_),
    .B(_17131_),
    .Y(_17134_));
 sky130_fd_sc_hd__nand3_4 _39505_ (.A(_17132_),
    .B(_17134_),
    .C(_16802_),
    .Y(_17135_));
 sky130_fd_sc_hd__a21o_1 _39506_ (.A1(_17128_),
    .A2(_17129_),
    .B1(_17130_),
    .X(_17136_));
 sky130_fd_sc_hd__nand2_1 _39507_ (.A(_17133_),
    .B(_17130_),
    .Y(_17137_));
 sky130_fd_sc_hd__nand3_2 _39508_ (.A(_17136_),
    .B(_17137_),
    .C(_16977_),
    .Y(_17138_));
 sky130_fd_sc_hd__nand3_2 _39509_ (.A(_17124_),
    .B(_17135_),
    .C(_17138_),
    .Y(_17139_));
 sky130_vsdinv _39510_ (.A(_17139_),
    .Y(_17140_));
 sky130_fd_sc_hd__nand2_1 _39511_ (.A(_17138_),
    .B(_17135_),
    .Y(_17141_));
 sky130_fd_sc_hd__a21oi_1 _39512_ (.A1(_16949_),
    .A2(_16952_),
    .B1(_17123_),
    .Y(_17142_));
 sky130_fd_sc_hd__nand2_1 _39513_ (.A(_17141_),
    .B(_17142_),
    .Y(_17143_));
 sky130_vsdinv _39514_ (.A(_16975_),
    .Y(_17144_));
 sky130_fd_sc_hd__a21oi_2 _39515_ (.A1(_16802_),
    .A2(_16976_),
    .B1(_17144_),
    .Y(_17145_));
 sky130_vsdinv _39516_ (.A(_17145_),
    .Y(_17146_));
 sky130_fd_sc_hd__nand2_2 _39517_ (.A(_17143_),
    .B(_17146_),
    .Y(_17147_));
 sky130_fd_sc_hd__nand2_1 _39518_ (.A(_17139_),
    .B(_17143_),
    .Y(_17148_));
 sky130_fd_sc_hd__nand2_2 _39519_ (.A(_17148_),
    .B(_17145_),
    .Y(_17149_));
 sky130_fd_sc_hd__o21a_1 _39520_ (.A1(_17140_),
    .A2(_17147_),
    .B1(_17149_),
    .X(_17150_));
 sky130_fd_sc_hd__o21ai_2 _39521_ (.A1(_17119_),
    .A2(_17122_),
    .B1(_17150_),
    .Y(_17151_));
 sky130_fd_sc_hd__a21o_1 _39522_ (.A1(_17115_),
    .A2(_17116_),
    .B1(_17118_),
    .X(_17152_));
 sky130_fd_sc_hd__nand3_4 _39523_ (.A(_17115_),
    .B(_17118_),
    .C(_17116_),
    .Y(_17153_));
 sky130_fd_sc_hd__o21ai_4 _39524_ (.A1(_17140_),
    .A2(_17147_),
    .B1(_17149_),
    .Y(_17154_));
 sky130_fd_sc_hd__nand3_2 _39525_ (.A(_17152_),
    .B(_17153_),
    .C(_17154_),
    .Y(_17155_));
 sky130_fd_sc_hd__nand3_4 _39526_ (.A(_17069_),
    .B(_17151_),
    .C(_17155_),
    .Y(_17156_));
 sky130_fd_sc_hd__o21ai_2 _39527_ (.A1(_17119_),
    .A2(_17122_),
    .B1(_17154_),
    .Y(_17157_));
 sky130_fd_sc_hd__o21ai_2 _39528_ (.A1(_16985_),
    .A2(_16963_),
    .B1(_16992_),
    .Y(_17158_));
 sky130_fd_sc_hd__nand3_2 _39529_ (.A(_17152_),
    .B(_17150_),
    .C(_17153_),
    .Y(_17159_));
 sky130_fd_sc_hd__nand3_4 _39530_ (.A(_17157_),
    .B(_17158_),
    .C(_17159_),
    .Y(_17160_));
 sky130_fd_sc_hd__nand2_1 _39531_ (.A(_17156_),
    .B(_17160_),
    .Y(_17161_));
 sky130_fd_sc_hd__nand2_2 _39532_ (.A(_16898_),
    .B(_16899_),
    .Y(_17162_));
 sky130_fd_sc_hd__a21o_2 _39533_ (.A1(_16787_),
    .A2(_16783_),
    .B1(_16709_),
    .X(_17163_));
 sky130_fd_sc_hd__nand2_1 _39534_ (.A(_17162_),
    .B(_17163_),
    .Y(_17164_));
 sky130_fd_sc_hd__or2_4 _39535_ (.A(_15753_),
    .B(_17164_),
    .X(_17165_));
 sky130_fd_sc_hd__nand2_2 _39536_ (.A(_17164_),
    .B(_15754_),
    .Y(_17166_));
 sky130_fd_sc_hd__nand2_4 _39537_ (.A(_17165_),
    .B(_17166_),
    .Y(_17167_));
 sky130_fd_sc_hd__a21o_2 _39538_ (.A1(_16984_),
    .A2(_16980_),
    .B1(_17167_),
    .X(_17168_));
 sky130_fd_sc_hd__nand3_4 _39539_ (.A(_17167_),
    .B(_16984_),
    .C(_16980_),
    .Y(_17169_));
 sky130_fd_sc_hd__nand2_2 _39540_ (.A(_16905_),
    .B(_17163_),
    .Y(_17170_));
 sky130_fd_sc_hd__a21oi_4 _39541_ (.A1(_17168_),
    .A2(_17169_),
    .B1(_17170_),
    .Y(_17171_));
 sky130_vsdinv _39542_ (.A(_17163_),
    .Y(_17172_));
 sky130_fd_sc_hd__o211a_1 _39543_ (.A1(_16906_),
    .A2(_17172_),
    .B1(_17169_),
    .C1(_17168_),
    .X(_17173_));
 sky130_fd_sc_hd__nor2_4 _39544_ (.A(_17171_),
    .B(_17173_),
    .Y(_17174_));
 sky130_fd_sc_hd__nand2_2 _39545_ (.A(_17161_),
    .B(_17174_),
    .Y(_17175_));
 sky130_fd_sc_hd__nand3b_4 _39546_ (.A_N(_17174_),
    .B(_17156_),
    .C(_17160_),
    .Y(_17176_));
 sky130_fd_sc_hd__o22ai_1 _39547_ (.A1(_16912_),
    .A2(_16914_),
    .B1(_16996_),
    .B2(_16999_),
    .Y(_17177_));
 sky130_fd_sc_hd__nand2_2 _39548_ (.A(_17177_),
    .B(_17004_),
    .Y(_17178_));
 sky130_fd_sc_hd__a21oi_4 _39549_ (.A1(_17175_),
    .A2(_17176_),
    .B1(_17178_),
    .Y(_17179_));
 sky130_fd_sc_hd__nand3_4 _39550_ (.A(_17175_),
    .B(_17178_),
    .C(_17176_),
    .Y(_17180_));
 sky130_fd_sc_hd__nand2_1 _39551_ (.A(_16913_),
    .B(_16908_),
    .Y(_17181_));
 sky130_fd_sc_hd__nand2_2 _39552_ (.A(_17181_),
    .B(_16147_),
    .Y(_17182_));
 sky130_fd_sc_hd__nand3_4 _39553_ (.A(_16149_),
    .B(_16908_),
    .C(_16913_),
    .Y(_17183_));
 sky130_fd_sc_hd__a21oi_4 _39554_ (.A1(_17182_),
    .A2(_17183_),
    .B1(_16484_),
    .Y(_17184_));
 sky130_fd_sc_hd__and3_1 _39555_ (.A(_17182_),
    .B(_17183_),
    .C(_16482_),
    .X(_17185_));
 sky130_fd_sc_hd__nor2_4 _39556_ (.A(_17184_),
    .B(_17185_),
    .Y(_17186_));
 sky130_fd_sc_hd__nand2_2 _39557_ (.A(_17180_),
    .B(_17186_),
    .Y(_17187_));
 sky130_fd_sc_hd__nand2_2 _39558_ (.A(_17022_),
    .B(_17023_),
    .Y(_17188_));
 sky130_fd_sc_hd__or2b_1 _39559_ (.A(_16912_),
    .B_N(_16913_),
    .X(_17189_));
 sky130_fd_sc_hd__o22ai_4 _39560_ (.A1(_16996_),
    .A2(_16999_),
    .B1(_17189_),
    .B2(_16995_),
    .Y(_17190_));
 sky130_fd_sc_hd__or2_1 _39561_ (.A(_17171_),
    .B(_17173_),
    .X(_17191_));
 sky130_fd_sc_hd__nand2_1 _39562_ (.A(_17161_),
    .B(_17191_),
    .Y(_17192_));
 sky130_fd_sc_hd__nand3_2 _39563_ (.A(_17156_),
    .B(_17160_),
    .C(_17174_),
    .Y(_17193_));
 sky130_fd_sc_hd__nand3_4 _39564_ (.A(_17190_),
    .B(_17192_),
    .C(_17193_),
    .Y(_17194_));
 sky130_fd_sc_hd__o2bb2ai_1 _39565_ (.A1_N(_17180_),
    .A2_N(_17194_),
    .B1(_17185_),
    .B2(_17184_),
    .Y(_17195_));
 sky130_fd_sc_hd__o2111ai_4 _39566_ (.A1(_17179_),
    .A2(_17187_),
    .B1(_17021_),
    .C1(_17188_),
    .D1(_17195_),
    .Y(_17196_));
 sky130_fd_sc_hd__a31oi_4 _39567_ (.A1(_17001_),
    .A2(_17006_),
    .A3(_17005_),
    .B1(_17017_),
    .Y(_17197_));
 sky130_fd_sc_hd__nand3b_4 _39568_ (.A_N(_17186_),
    .B(_17194_),
    .C(_17180_),
    .Y(_17198_));
 sky130_fd_sc_hd__nand2_1 _39569_ (.A(_17194_),
    .B(_17180_),
    .Y(_17199_));
 sky130_fd_sc_hd__nand2_4 _39570_ (.A(_17199_),
    .B(_17186_),
    .Y(_17200_));
 sky130_fd_sc_hd__o211ai_4 _39571_ (.A1(_17007_),
    .A2(_17197_),
    .B1(_17198_),
    .C1(_17200_),
    .Y(_17201_));
 sky130_vsdinv _39572_ (.A(_17011_),
    .Y(_17202_));
 sky130_fd_sc_hd__clkbuf_4 _39573_ (.A(_16482_),
    .X(_17203_));
 sky130_fd_sc_hd__a21oi_4 _39574_ (.A1(_17202_),
    .A2(_17203_),
    .B1(_17015_),
    .Y(_17204_));
 sky130_fd_sc_hd__nor2_4 _39575_ (.A(_14903_),
    .B(_17204_),
    .Y(_17205_));
 sky130_fd_sc_hd__a21o_1 _39576_ (.A1(_17202_),
    .A2(_17203_),
    .B1(_17015_),
    .X(_17206_));
 sky130_fd_sc_hd__nor2_4 _39577_ (.A(_14329_),
    .B(_17206_),
    .Y(_17207_));
 sky130_fd_sc_hd__nor2_4 _39578_ (.A(_17205_),
    .B(_17207_),
    .Y(_17208_));
 sky130_vsdinv _39579_ (.A(_17208_),
    .Y(_17209_));
 sky130_fd_sc_hd__nand3_2 _39580_ (.A(_17196_),
    .B(_17201_),
    .C(_17209_),
    .Y(_17210_));
 sky130_fd_sc_hd__a21o_1 _39581_ (.A1(_17196_),
    .A2(_17201_),
    .B1(_17209_),
    .X(_17211_));
 sky130_fd_sc_hd__o211ai_4 _39582_ (.A1(_17067_),
    .A2(_17068_),
    .B1(_17210_),
    .C1(_17211_),
    .Y(_17212_));
 sky130_fd_sc_hd__nand2_1 _39583_ (.A(_17026_),
    .B(_17028_),
    .Y(_17213_));
 sky130_fd_sc_hd__nand3_4 _39584_ (.A(_17196_),
    .B(_17201_),
    .C(_17208_),
    .Y(_17214_));
 sky130_fd_sc_hd__nand2_1 _39585_ (.A(_17025_),
    .B(_17043_),
    .Y(_17215_));
 sky130_fd_sc_hd__o2bb2ai_4 _39586_ (.A1_N(_17201_),
    .A2_N(_17196_),
    .B1(_17207_),
    .B2(_17205_),
    .Y(_17216_));
 sky130_fd_sc_hd__o2111ai_4 _39587_ (.A1(_17020_),
    .A2(_17213_),
    .B1(_17214_),
    .C1(_17215_),
    .D1(_17216_),
    .Y(_17217_));
 sky130_fd_sc_hd__a21oi_1 _39588_ (.A1(_17212_),
    .A2(_17217_),
    .B1(_17042_),
    .Y(_17218_));
 sky130_fd_sc_hd__and3_1 _39589_ (.A(_17212_),
    .B(_17217_),
    .C(_17042_),
    .X(_17219_));
 sky130_vsdinv _39590_ (.A(_17044_),
    .Y(_17220_));
 sky130_fd_sc_hd__nand2_1 _39591_ (.A(_17037_),
    .B(_17039_),
    .Y(_17221_));
 sky130_fd_sc_hd__o2bb2ai_2 _39592_ (.A1_N(_16864_),
    .A2_N(_17049_),
    .B1(_17220_),
    .B2(_17221_),
    .Y(_17222_));
 sky130_fd_sc_hd__o21bai_2 _39593_ (.A1(_17218_),
    .A2(_17219_),
    .B1_N(_17222_),
    .Y(_17223_));
 sky130_fd_sc_hd__a21o_1 _39594_ (.A1(_17212_),
    .A2(_17217_),
    .B1(_17042_),
    .X(_17224_));
 sky130_fd_sc_hd__a21oi_4 _39595_ (.A1(_17025_),
    .A2(_17043_),
    .B1(_17067_),
    .Y(_17225_));
 sky130_fd_sc_hd__a31oi_4 _39596_ (.A1(_17225_),
    .A2(_17214_),
    .A3(_17216_),
    .B1(_17041_),
    .Y(_17226_));
 sky130_fd_sc_hd__nand2_1 _39597_ (.A(_17226_),
    .B(_17212_),
    .Y(_17227_));
 sky130_fd_sc_hd__nand3_4 _39598_ (.A(_17224_),
    .B(_17227_),
    .C(_17222_),
    .Y(_17228_));
 sky130_fd_sc_hd__nand2_1 _39599_ (.A(_17223_),
    .B(_17228_),
    .Y(_17229_));
 sky130_fd_sc_hd__a21oi_2 _39600_ (.A1(_17064_),
    .A2(_17066_),
    .B1(_17229_),
    .Y(_17230_));
 sky130_fd_sc_hd__and3_1 _39601_ (.A(_17064_),
    .B(_17229_),
    .C(_17066_),
    .X(_17231_));
 sky130_fd_sc_hd__nor2_1 _39602_ (.A(_17230_),
    .B(_17231_),
    .Y(_02673_));
 sky130_fd_sc_hd__nand2_2 _39603_ (.A(_17188_),
    .B(_17021_),
    .Y(_17232_));
 sky130_fd_sc_hd__a21oi_4 _39604_ (.A1(_17200_),
    .A2(_17198_),
    .B1(_17232_),
    .Y(_17233_));
 sky130_fd_sc_hd__a21oi_2 _39605_ (.A1(_17201_),
    .A2(_17209_),
    .B1(_17233_),
    .Y(_17234_));
 sky130_fd_sc_hd__nand2_1 _39606_ (.A(_17147_),
    .B(_17139_),
    .Y(_17235_));
 sky130_fd_sc_hd__a21o_2 _39607_ (.A1(_17166_),
    .A2(_17165_),
    .B1(_17235_),
    .X(_17236_));
 sky130_fd_sc_hd__and2_2 _39608_ (.A(_17165_),
    .B(_17166_),
    .X(_17237_));
 sky130_fd_sc_hd__nand2_2 _39609_ (.A(_17237_),
    .B(_17235_),
    .Y(_17238_));
 sky130_fd_sc_hd__nand2_4 _39610_ (.A(_17165_),
    .B(_17163_),
    .Y(_17239_));
 sky130_fd_sc_hd__a21oi_4 _39611_ (.A1(_17236_),
    .A2(_17238_),
    .B1(_17239_),
    .Y(_17240_));
 sky130_fd_sc_hd__nand3_1 _39612_ (.A(_17236_),
    .B(_17238_),
    .C(_17239_),
    .Y(_17241_));
 sky130_vsdinv _39613_ (.A(_17241_),
    .Y(_17242_));
 sky130_vsdinv _39614_ (.A(_19613_),
    .Y(_17243_));
 sky130_vsdinv _39615_ (.A(_19609_),
    .Y(_17244_));
 sky130_fd_sc_hd__clkbuf_2 _39616_ (.A(_13007_),
    .X(_17245_));
 sky130_fd_sc_hd__a21oi_2 _39617_ (.A1(_19613_),
    .A2(_19619_),
    .B1(_17245_),
    .Y(_17246_));
 sky130_fd_sc_hd__a211o_1 _39618_ (.A1(_17243_),
    .A2(_07833_),
    .B1(_17244_),
    .C1(_17246_),
    .X(_17247_));
 sky130_fd_sc_hd__a31o_1 _39619_ (.A1(_17244_),
    .A2(_17243_),
    .A3(_07833_),
    .B1(net465),
    .X(_17248_));
 sky130_vsdinv _39620_ (.A(_17248_),
    .Y(_17249_));
 sky130_fd_sc_hd__nand2_1 _39621_ (.A(_17247_),
    .B(_17249_),
    .Y(_17250_));
 sky130_fd_sc_hd__nor2_1 _39622_ (.A(_17250_),
    .B(_16977_),
    .Y(_17251_));
 sky130_vsdinv _39623_ (.A(_17251_),
    .Y(_17252_));
 sky130_fd_sc_hd__nand2_2 _39624_ (.A(_16977_),
    .B(_17250_),
    .Y(_17253_));
 sky130_fd_sc_hd__a21oi_2 _39625_ (.A1(_17105_),
    .A2(_17106_),
    .B1(_17107_),
    .Y(_17254_));
 sky130_fd_sc_hd__o21ai_4 _39626_ (.A1(_17111_),
    .A2(_17254_),
    .B1(_17109_),
    .Y(_17255_));
 sky130_fd_sc_hd__a21o_1 _39627_ (.A1(_17252_),
    .A2(_17253_),
    .B1(_17255_),
    .X(_17256_));
 sky130_fd_sc_hd__nand3_4 _39628_ (.A(_17255_),
    .B(_17253_),
    .C(_17252_),
    .Y(_17257_));
 sky130_fd_sc_hd__nand2_2 _39629_ (.A(_17135_),
    .B(_17132_),
    .Y(_17258_));
 sky130_fd_sc_hd__a21oi_4 _39630_ (.A1(_17256_),
    .A2(_17257_),
    .B1(_17258_),
    .Y(_17259_));
 sky130_vsdinv _39631_ (.A(_17258_),
    .Y(_17260_));
 sky130_fd_sc_hd__nand2_2 _39632_ (.A(_17256_),
    .B(_17257_),
    .Y(_17261_));
 sky130_fd_sc_hd__nor2_4 _39633_ (.A(_17260_),
    .B(_17261_),
    .Y(_17262_));
 sky130_fd_sc_hd__o311a_2 _39634_ (.A1(_17074_),
    .A2(_17075_),
    .A3(_17077_),
    .B1(_17086_),
    .C1(_17085_),
    .X(_17263_));
 sky130_fd_sc_hd__nand2_1 _39635_ (.A(_15806_),
    .B(_19841_),
    .Y(_17264_));
 sky130_fd_sc_hd__o22a_1 _39636_ (.A1(_16159_),
    .A2(_10617_),
    .B1(_15932_),
    .B2(_10497_),
    .X(_17265_));
 sky130_fd_sc_hd__a31o_1 _39637_ (.A1(_19845_),
    .A2(_19850_),
    .A3(_15930_),
    .B1(_17265_),
    .X(_17266_));
 sky130_fd_sc_hd__nor2_2 _39638_ (.A(_17264_),
    .B(_17266_),
    .Y(_17267_));
 sky130_fd_sc_hd__and2_1 _39639_ (.A(_17266_),
    .B(_17264_),
    .X(_17268_));
 sky130_fd_sc_hd__nor2_4 _39640_ (.A(_17267_),
    .B(_17268_),
    .Y(_17269_));
 sky130_fd_sc_hd__nand2_2 _39641_ (.A(_19580_),
    .B(_19853_),
    .Y(_17270_));
 sky130_fd_sc_hd__and4_2 _39642_ (.A(_10466_),
    .B(_15937_),
    .C(_15821_),
    .D(_14501_),
    .X(_17271_));
 sky130_fd_sc_hd__o22a_2 _39643_ (.A1(_19860_),
    .A2(_16352_),
    .B1(_15817_),
    .B2(_09929_),
    .X(_17272_));
 sky130_fd_sc_hd__or3_4 _39644_ (.A(_17270_),
    .B(_17271_),
    .C(_17272_),
    .X(_17273_));
 sky130_fd_sc_hd__o21ai_4 _39645_ (.A1(_17271_),
    .A2(_17272_),
    .B1(_17270_),
    .Y(_17274_));
 sky130_fd_sc_hd__nor2_4 _39646_ (.A(_17071_),
    .B(_17072_),
    .Y(_17275_));
 sky130_fd_sc_hd__o2bb2ai_4 _39647_ (.A1_N(_17273_),
    .A2_N(_17274_),
    .B1(_17073_),
    .B2(_17275_),
    .Y(_17276_));
 sky130_fd_sc_hd__nor2_2 _39648_ (.A(_17073_),
    .B(_17275_),
    .Y(_17277_));
 sky130_fd_sc_hd__nand3_4 _39649_ (.A(_17273_),
    .B(_17274_),
    .C(_17277_),
    .Y(_17278_));
 sky130_fd_sc_hd__nand3_4 _39650_ (.A(_17269_),
    .B(_17276_),
    .C(_17278_),
    .Y(_17279_));
 sky130_fd_sc_hd__a21o_1 _39651_ (.A1(_17276_),
    .A2(_17278_),
    .B1(_17269_),
    .X(_17280_));
 sky130_fd_sc_hd__o211ai_4 _39652_ (.A1(_17078_),
    .A2(_17263_),
    .B1(_17279_),
    .C1(_17280_),
    .Y(_17281_));
 sky130_fd_sc_hd__a21oi_2 _39653_ (.A1(_17276_),
    .A2(_17278_),
    .B1(_17269_),
    .Y(_17282_));
 sky130_fd_sc_hd__a21oi_1 _39654_ (.A1(_19594_),
    .A2(_19842_),
    .B1(_17266_),
    .Y(_17283_));
 sky130_fd_sc_hd__and3_1 _39655_ (.A(_17266_),
    .B(_19594_),
    .C(_19842_),
    .X(_17284_));
 sky130_fd_sc_hd__o211a_1 _39656_ (.A1(_17283_),
    .A2(_17284_),
    .B1(_17278_),
    .C1(_17276_),
    .X(_17285_));
 sky130_fd_sc_hd__nor2_2 _39657_ (.A(_17078_),
    .B(_17263_),
    .Y(_17286_));
 sky130_fd_sc_hd__o21ai_4 _39658_ (.A1(_17282_),
    .A2(_17285_),
    .B1(_17286_),
    .Y(_17287_));
 sky130_fd_sc_hd__clkbuf_2 _39659_ (.A(_13309_),
    .X(_17288_));
 sky130_fd_sc_hd__nor2_1 _39660_ (.A(_16940_),
    .B(_15780_),
    .Y(_17289_));
 sky130_fd_sc_hd__or3_4 _39661_ (.A(_16184_),
    .B(_17288_),
    .C(_17289_),
    .X(_17290_));
 sky130_fd_sc_hd__o21ai_2 _39662_ (.A1(_16184_),
    .A2(_17288_),
    .B1(_17289_),
    .Y(_17291_));
 sky130_fd_sc_hd__nand2_2 _39663_ (.A(_19605_),
    .B(_19828_),
    .Y(_17292_));
 sky130_fd_sc_hd__a21o_1 _39664_ (.A1(_17290_),
    .A2(_17291_),
    .B1(_17292_),
    .X(_17293_));
 sky130_fd_sc_hd__nand3_4 _39665_ (.A(_17290_),
    .B(_17291_),
    .C(_17292_),
    .Y(_17294_));
 sky130_fd_sc_hd__a21o_1 _39666_ (.A1(_17084_),
    .A2(_17081_),
    .B1(_17083_),
    .X(_17295_));
 sky130_fd_sc_hd__a21o_2 _39667_ (.A1(_17293_),
    .A2(_17294_),
    .B1(_17295_),
    .X(_17296_));
 sky130_fd_sc_hd__nand3_4 _39668_ (.A(_17293_),
    .B(_17295_),
    .C(_17294_),
    .Y(_17297_));
 sky130_fd_sc_hd__a21o_2 _39669_ (.A1(_17104_),
    .A2(_17099_),
    .B1(_17102_),
    .X(_17298_));
 sky130_fd_sc_hd__and3_1 _39670_ (.A(_17296_),
    .B(_17297_),
    .C(_17298_),
    .X(_17299_));
 sky130_fd_sc_hd__a21oi_2 _39671_ (.A1(_17296_),
    .A2(_17297_),
    .B1(_17298_),
    .Y(_17300_));
 sky130_fd_sc_hd__o2bb2ai_4 _39672_ (.A1_N(_17281_),
    .A2_N(_17287_),
    .B1(_17299_),
    .B2(_17300_),
    .Y(_17301_));
 sky130_fd_sc_hd__nand2_1 _39673_ (.A(_17296_),
    .B(_17297_),
    .Y(_17302_));
 sky130_fd_sc_hd__nand2_1 _39674_ (.A(_17302_),
    .B(_17298_),
    .Y(_17303_));
 sky130_fd_sc_hd__nand3b_1 _39675_ (.A_N(_17298_),
    .B(_17296_),
    .C(_17297_),
    .Y(_17304_));
 sky130_fd_sc_hd__nand2_1 _39676_ (.A(_17303_),
    .B(_17304_),
    .Y(_17305_));
 sky130_fd_sc_hd__nand3_4 _39677_ (.A(_17305_),
    .B(_17281_),
    .C(_17287_),
    .Y(_17306_));
 sky130_fd_sc_hd__nand2_2 _39678_ (.A(_17121_),
    .B(_17094_),
    .Y(_17307_));
 sky130_fd_sc_hd__a21oi_2 _39679_ (.A1(_17301_),
    .A2(_17306_),
    .B1(_17307_),
    .Y(_17308_));
 sky130_fd_sc_hd__nand2_1 _39680_ (.A(_17096_),
    .B(_17097_),
    .Y(_17309_));
 sky130_fd_sc_hd__o21a_1 _39681_ (.A1(_17070_),
    .A2(_17309_),
    .B1(_17114_),
    .X(_17310_));
 sky130_fd_sc_hd__o211a_2 _39682_ (.A1(_17120_),
    .A2(_17310_),
    .B1(_17306_),
    .C1(_17301_),
    .X(_17311_));
 sky130_fd_sc_hd__o22ai_4 _39683_ (.A1(_17259_),
    .A2(_17262_),
    .B1(_17308_),
    .B2(_17311_),
    .Y(_17312_));
 sky130_fd_sc_hd__a21o_1 _39684_ (.A1(_17301_),
    .A2(_17306_),
    .B1(_17307_),
    .X(_17313_));
 sky130_fd_sc_hd__nand3_2 _39685_ (.A(_17301_),
    .B(_17306_),
    .C(_17307_),
    .Y(_17314_));
 sky130_fd_sc_hd__nor2_4 _39686_ (.A(_17259_),
    .B(_17262_),
    .Y(_17315_));
 sky130_fd_sc_hd__nand3_4 _39687_ (.A(_17313_),
    .B(_17314_),
    .C(_17315_),
    .Y(_17316_));
 sky130_fd_sc_hd__o21ai_4 _39688_ (.A1(_17154_),
    .A2(_17119_),
    .B1(_17153_),
    .Y(_17317_));
 sky130_fd_sc_hd__a21oi_4 _39689_ (.A1(_17312_),
    .A2(_17316_),
    .B1(_17317_),
    .Y(_17318_));
 sky130_fd_sc_hd__nor2_1 _39690_ (.A(_17154_),
    .B(_17119_),
    .Y(_17319_));
 sky130_fd_sc_hd__o211a_1 _39691_ (.A1(_17122_),
    .A2(_17319_),
    .B1(_17316_),
    .C1(_17312_),
    .X(_17320_));
 sky130_fd_sc_hd__o22ai_4 _39692_ (.A1(_17240_),
    .A2(_17242_),
    .B1(_17318_),
    .B2(_17320_),
    .Y(_17321_));
 sky130_fd_sc_hd__nand2_1 _39693_ (.A(_17156_),
    .B(_17174_),
    .Y(_17322_));
 sky130_fd_sc_hd__nand2_1 _39694_ (.A(_17322_),
    .B(_17160_),
    .Y(_17323_));
 sky130_fd_sc_hd__a21o_1 _39695_ (.A1(_17312_),
    .A2(_17316_),
    .B1(_17317_),
    .X(_17324_));
 sky130_fd_sc_hd__nand3_4 _39696_ (.A(_17312_),
    .B(_17317_),
    .C(_17316_),
    .Y(_17325_));
 sky130_fd_sc_hd__and2_1 _39697_ (.A(_17238_),
    .B(_17239_),
    .X(_17326_));
 sky130_fd_sc_hd__a21oi_2 _39698_ (.A1(_17326_),
    .A2(_17236_),
    .B1(_17240_),
    .Y(_17327_));
 sky130_fd_sc_hd__nand3_2 _39699_ (.A(_17324_),
    .B(_17325_),
    .C(_17327_),
    .Y(_17328_));
 sky130_fd_sc_hd__nand3_4 _39700_ (.A(_17321_),
    .B(_17323_),
    .C(_17328_),
    .Y(_17329_));
 sky130_fd_sc_hd__o21ai_2 _39701_ (.A1(_17318_),
    .A2(_17320_),
    .B1(_17327_),
    .Y(_17330_));
 sky130_fd_sc_hd__a21boi_2 _39702_ (.A1(_17156_),
    .A2(_17174_),
    .B1_N(_17160_),
    .Y(_17331_));
 sky130_fd_sc_hd__a21o_1 _39703_ (.A1(_17236_),
    .A2(_17326_),
    .B1(_17240_),
    .X(_17332_));
 sky130_fd_sc_hd__nand3_2 _39704_ (.A(_17324_),
    .B(_17332_),
    .C(_17325_),
    .Y(_17333_));
 sky130_fd_sc_hd__nand3_4 _39705_ (.A(_17330_),
    .B(_17331_),
    .C(_17333_),
    .Y(_17334_));
 sky130_fd_sc_hd__nand3_2 _39706_ (.A(_17168_),
    .B(_17170_),
    .C(_17169_),
    .Y(_17335_));
 sky130_fd_sc_hd__a21o_1 _39707_ (.A1(_17335_),
    .A2(_17168_),
    .B1(_16149_),
    .X(_17336_));
 sky130_fd_sc_hd__nand3_2 _39708_ (.A(_16149_),
    .B(_17335_),
    .C(_17168_),
    .Y(_17337_));
 sky130_fd_sc_hd__and3_1 _39709_ (.A(_17336_),
    .B(_16482_),
    .C(_17337_),
    .X(_17338_));
 sky130_fd_sc_hd__a21oi_2 _39710_ (.A1(_17336_),
    .A2(_17337_),
    .B1(_16484_),
    .Y(_17339_));
 sky130_fd_sc_hd__o2bb2ai_2 _39711_ (.A1_N(_17329_),
    .A2_N(_17334_),
    .B1(_17338_),
    .B2(_17339_),
    .Y(_17340_));
 sky130_fd_sc_hd__nand2_1 _39712_ (.A(_17187_),
    .B(_17194_),
    .Y(_17341_));
 sky130_fd_sc_hd__nor2_2 _39713_ (.A(_17339_),
    .B(_17338_),
    .Y(_17342_));
 sky130_fd_sc_hd__nand3_2 _39714_ (.A(_17334_),
    .B(_17329_),
    .C(_17342_),
    .Y(_17343_));
 sky130_fd_sc_hd__nand3_4 _39715_ (.A(_17340_),
    .B(_17341_),
    .C(_17343_),
    .Y(_17344_));
 sky130_fd_sc_hd__nand2_1 _39716_ (.A(_17334_),
    .B(_17329_),
    .Y(_17345_));
 sky130_fd_sc_hd__nand2_1 _39717_ (.A(_17345_),
    .B(_17342_),
    .Y(_17346_));
 sky130_fd_sc_hd__a21oi_2 _39718_ (.A1(_17180_),
    .A2(_17186_),
    .B1(_17179_),
    .Y(_17347_));
 sky130_fd_sc_hd__nand3b_2 _39719_ (.A_N(_17342_),
    .B(_17334_),
    .C(_17329_),
    .Y(_17348_));
 sky130_fd_sc_hd__nand3_4 _39720_ (.A(_17346_),
    .B(_17347_),
    .C(_17348_),
    .Y(_17349_));
 sky130_fd_sc_hd__nand2_1 _39721_ (.A(_17183_),
    .B(_17203_),
    .Y(_17350_));
 sky130_fd_sc_hd__nand2_2 _39722_ (.A(_17350_),
    .B(_17182_),
    .Y(_17351_));
 sky130_fd_sc_hd__nor2_1 _39723_ (.A(_14331_),
    .B(_17351_),
    .Y(_17352_));
 sky130_fd_sc_hd__buf_4 _39724_ (.A(_16675_),
    .X(_17353_));
 sky130_vsdinv _39725_ (.A(_17351_),
    .Y(_17354_));
 sky130_fd_sc_hd__nor2_1 _39726_ (.A(_17353_),
    .B(_17354_),
    .Y(_17355_));
 sky130_fd_sc_hd__o2bb2ai_2 _39727_ (.A1_N(_17344_),
    .A2_N(_17349_),
    .B1(_17352_),
    .B2(_17355_),
    .Y(_17356_));
 sky130_fd_sc_hd__nor2_2 _39728_ (.A(_16317_),
    .B(_17351_),
    .Y(_17357_));
 sky130_fd_sc_hd__nor2_1 _39729_ (.A(_14330_),
    .B(_17354_),
    .Y(_17358_));
 sky130_fd_sc_hd__nor2_2 _39730_ (.A(_17357_),
    .B(_17358_),
    .Y(_17359_));
 sky130_fd_sc_hd__nand3b_2 _39731_ (.A_N(_17359_),
    .B(_17349_),
    .C(_17344_),
    .Y(_17360_));
 sky130_fd_sc_hd__nand3_4 _39732_ (.A(_17234_),
    .B(_17356_),
    .C(_17360_),
    .Y(_17361_));
 sky130_fd_sc_hd__a31oi_4 _39733_ (.A1(_17232_),
    .A2(_17200_),
    .A3(_17198_),
    .B1(_17208_),
    .Y(_17362_));
 sky130_fd_sc_hd__nand3_2 _39734_ (.A(_17349_),
    .B(_17344_),
    .C(_17359_),
    .Y(_17363_));
 sky130_fd_sc_hd__buf_2 _39735_ (.A(_17358_),
    .X(_17364_));
 sky130_fd_sc_hd__o2bb2ai_2 _39736_ (.A1_N(_17344_),
    .A2_N(_17349_),
    .B1(_17364_),
    .B2(_17357_),
    .Y(_17365_));
 sky130_fd_sc_hd__o211ai_4 _39737_ (.A1(_17233_),
    .A2(_17362_),
    .B1(_17363_),
    .C1(_17365_),
    .Y(_17366_));
 sky130_fd_sc_hd__nor2_2 _39738_ (.A(net410),
    .B(_17204_),
    .Y(_17367_));
 sky130_fd_sc_hd__and3_4 _39739_ (.A(_17361_),
    .B(_17366_),
    .C(_17367_),
    .X(_17368_));
 sky130_vsdinv _39740_ (.A(_17367_),
    .Y(_17369_));
 sky130_fd_sc_hd__nand2_2 _39741_ (.A(_17361_),
    .B(_17366_),
    .Y(_17370_));
 sky130_fd_sc_hd__a21oi_4 _39742_ (.A1(_17214_),
    .A2(_17216_),
    .B1(_17225_),
    .Y(_17371_));
 sky130_fd_sc_hd__o2bb2ai_4 _39743_ (.A1_N(_17369_),
    .A2_N(_17370_),
    .B1(_17371_),
    .B2(_17226_),
    .Y(_17372_));
 sky130_fd_sc_hd__a21oi_2 _39744_ (.A1(_17361_),
    .A2(_17366_),
    .B1(_17367_),
    .Y(_17373_));
 sky130_fd_sc_hd__nor2_2 _39745_ (.A(_17371_),
    .B(_17226_),
    .Y(_17374_));
 sky130_fd_sc_hd__o21ai_4 _39746_ (.A1(_17373_),
    .A2(_17368_),
    .B1(_17374_),
    .Y(_17375_));
 sky130_fd_sc_hd__o21a_1 _39747_ (.A1(_17368_),
    .A2(_17372_),
    .B1(_17375_),
    .X(_17376_));
 sky130_fd_sc_hd__nand3b_1 _39748_ (.A_N(_17230_),
    .B(_17228_),
    .C(_17376_),
    .Y(_17377_));
 sky130_vsdinv _39749_ (.A(_17228_),
    .Y(_17378_));
 sky130_fd_sc_hd__o21bai_1 _39750_ (.A1(_17378_),
    .A2(_17230_),
    .B1_N(_17376_),
    .Y(_17379_));
 sky130_fd_sc_hd__nand2_1 _39751_ (.A(_17377_),
    .B(_17379_),
    .Y(_02674_));
 sky130_fd_sc_hd__o21ai_4 _39752_ (.A1(_17318_),
    .A2(_17332_),
    .B1(_17325_),
    .Y(_17380_));
 sky130_fd_sc_hd__nand2_2 _39753_ (.A(_17279_),
    .B(_17278_),
    .Y(_17381_));
 sky130_fd_sc_hd__nand2_1 _39754_ (.A(_19581_),
    .B(_19850_),
    .Y(_17382_));
 sky130_fd_sc_hd__or4_4 _39755_ (.A(_19856_),
    .B(_16352_),
    .C(_15817_),
    .D(_13855_),
    .X(_17383_));
 sky130_fd_sc_hd__a22o_1 _39756_ (.A1(_19578_),
    .A2(_19853_),
    .B1(_09929_),
    .B2(_11293_),
    .X(_17384_));
 sky130_fd_sc_hd__nand2_1 _39757_ (.A(_17383_),
    .B(_17384_),
    .Y(_17385_));
 sky130_fd_sc_hd__or2_4 _39758_ (.A(_17382_),
    .B(_17385_),
    .X(_17386_));
 sky130_fd_sc_hd__nand2_2 _39759_ (.A(_17385_),
    .B(_17382_),
    .Y(_17387_));
 sky130_fd_sc_hd__nand2_1 _39760_ (.A(_17386_),
    .B(_17387_),
    .Y(_17388_));
 sky130_vsdinv _39761_ (.A(_17271_),
    .Y(_17389_));
 sky130_fd_sc_hd__nand2_2 _39762_ (.A(_17273_),
    .B(_17389_),
    .Y(_17390_));
 sky130_vsdinv _39763_ (.A(_17390_),
    .Y(_17391_));
 sky130_fd_sc_hd__nand2_2 _39764_ (.A(_17388_),
    .B(_17391_),
    .Y(_17392_));
 sky130_fd_sc_hd__nand3_4 _39765_ (.A(_17386_),
    .B(_17390_),
    .C(_17387_),
    .Y(_17393_));
 sky130_fd_sc_hd__nand2_1 _39766_ (.A(_15806_),
    .B(_19836_),
    .Y(_17394_));
 sky130_fd_sc_hd__nand2_2 _39767_ (.A(_19584_),
    .B(_19840_),
    .Y(_17395_));
 sky130_fd_sc_hd__a22o_1 _39768_ (.A1(_19584_),
    .A2(_19844_),
    .B1(_19588_),
    .B2(_10601_),
    .X(_17396_));
 sky130_fd_sc_hd__o31ai_4 _39769_ (.A1(_17395_),
    .A2(_15834_),
    .A3(_13900_),
    .B1(_17396_),
    .Y(_17397_));
 sky130_fd_sc_hd__nor2_1 _39770_ (.A(_17394_),
    .B(_17397_),
    .Y(_17398_));
 sky130_fd_sc_hd__and2_1 _39771_ (.A(_17397_),
    .B(_17394_),
    .X(_17399_));
 sky130_fd_sc_hd__or2_4 _39772_ (.A(_17398_),
    .B(_17399_),
    .X(_17400_));
 sky130_fd_sc_hd__nand3_2 _39773_ (.A(_17392_),
    .B(_17393_),
    .C(_17400_),
    .Y(_17401_));
 sky130_fd_sc_hd__nand2_1 _39774_ (.A(_17388_),
    .B(_17390_),
    .Y(_17402_));
 sky130_fd_sc_hd__nand3_2 _39775_ (.A(_17386_),
    .B(_17391_),
    .C(_17387_),
    .Y(_17403_));
 sky130_vsdinv _39776_ (.A(_17400_),
    .Y(_17404_));
 sky130_fd_sc_hd__nand3_2 _39777_ (.A(_17402_),
    .B(_17403_),
    .C(_17404_),
    .Y(_17405_));
 sky130_fd_sc_hd__nand3b_4 _39778_ (.A_N(_17381_),
    .B(_17401_),
    .C(_17405_),
    .Y(_17406_));
 sky130_fd_sc_hd__nand3_2 _39779_ (.A(_17392_),
    .B(_17393_),
    .C(_17404_),
    .Y(_17407_));
 sky130_fd_sc_hd__nand3_2 _39780_ (.A(_17402_),
    .B(_17403_),
    .C(_17400_),
    .Y(_17408_));
 sky130_fd_sc_hd__nand3_4 _39781_ (.A(_17407_),
    .B(_17408_),
    .C(_17381_),
    .Y(_17409_));
 sky130_fd_sc_hd__nand2_4 _39782_ (.A(_14218_),
    .B(_19604_),
    .Y(_17410_));
 sky130_fd_sc_hd__or4_4 _39783_ (.A(_16940_),
    .B(_16184_),
    .C(_13007_),
    .D(_13309_),
    .X(_17411_));
 sky130_fd_sc_hd__a22o_1 _39784_ (.A1(_19598_),
    .A2(_19831_),
    .B1(_19601_),
    .B2(_19827_),
    .X(_17412_));
 sky130_fd_sc_hd__nand2_1 _39785_ (.A(_17411_),
    .B(_17412_),
    .Y(_17413_));
 sky130_fd_sc_hd__or2_4 _39786_ (.A(_17410_),
    .B(_17413_),
    .X(_17414_));
 sky130_fd_sc_hd__nand2_2 _39787_ (.A(_17413_),
    .B(_17410_),
    .Y(_17415_));
 sky130_fd_sc_hd__a31o_2 _39788_ (.A1(_19846_),
    .A2(_19850_),
    .A3(_16946_),
    .B1(_17267_),
    .X(_17416_));
 sky130_fd_sc_hd__a21oi_4 _39789_ (.A1(_17414_),
    .A2(_17415_),
    .B1(_17416_),
    .Y(_17417_));
 sky130_fd_sc_hd__and3_1 _39790_ (.A(_17416_),
    .B(_17414_),
    .C(_17415_),
    .X(_17418_));
 sky130_fd_sc_hd__or4_4 _39791_ (.A(_16940_),
    .B(_16184_),
    .C(_17288_),
    .D(_15780_),
    .X(_17419_));
 sky130_fd_sc_hd__nand2_1 _39792_ (.A(_17293_),
    .B(_17419_),
    .Y(_17420_));
 sky130_fd_sc_hd__o21ai_1 _39793_ (.A1(_17417_),
    .A2(_17418_),
    .B1(_17420_),
    .Y(_17421_));
 sky130_vsdinv _39794_ (.A(_17420_),
    .Y(_17422_));
 sky130_fd_sc_hd__nand3_4 _39795_ (.A(_17416_),
    .B(_17414_),
    .C(_17415_),
    .Y(_17423_));
 sky130_fd_sc_hd__nand3b_1 _39796_ (.A_N(_17417_),
    .B(_17422_),
    .C(_17423_),
    .Y(_17424_));
 sky130_fd_sc_hd__nand2_2 _39797_ (.A(_17421_),
    .B(_17424_),
    .Y(_17425_));
 sky130_fd_sc_hd__a21o_2 _39798_ (.A1(_17406_),
    .A2(_17409_),
    .B1(_17425_),
    .X(_17426_));
 sky130_fd_sc_hd__nand3_4 _39799_ (.A(_17425_),
    .B(_17406_),
    .C(_17409_),
    .Y(_17427_));
 sky130_fd_sc_hd__nand2_2 _39800_ (.A(_17306_),
    .B(_17281_),
    .Y(_17428_));
 sky130_fd_sc_hd__a21oi_4 _39801_ (.A1(_17426_),
    .A2(_17427_),
    .B1(_17428_),
    .Y(_17429_));
 sky130_fd_sc_hd__and3_2 _39802_ (.A(_17426_),
    .B(_17428_),
    .C(_17427_),
    .X(_17430_));
 sky130_fd_sc_hd__nand2_2 _39803_ (.A(_17296_),
    .B(_17298_),
    .Y(_17431_));
 sky130_fd_sc_hd__or3_1 _39804_ (.A(_17126_),
    .B(_17244_),
    .C(_07833_),
    .X(_17432_));
 sky130_vsdinv _39805_ (.A(_17432_),
    .Y(_17433_));
 sky130_fd_sc_hd__nand2_4 _39806_ (.A(_16802_),
    .B(_17433_),
    .Y(_17434_));
 sky130_fd_sc_hd__a31o_1 _39807_ (.A1(_16787_),
    .A2(_16788_),
    .A3(_17249_),
    .B1(_17433_),
    .X(_17435_));
 sky130_fd_sc_hd__nor2_8 _39808_ (.A(_17249_),
    .B(_16802_),
    .Y(_17436_));
 sky130_fd_sc_hd__a21o_1 _39809_ (.A1(_17434_),
    .A2(_17435_),
    .B1(_17436_),
    .X(_17437_));
 sky130_fd_sc_hd__a21o_1 _39810_ (.A1(_17297_),
    .A2(_17431_),
    .B1(_17437_),
    .X(_17438_));
 sky130_fd_sc_hd__nand3_4 _39811_ (.A(_17437_),
    .B(_17297_),
    .C(_17431_),
    .Y(_17439_));
 sky130_fd_sc_hd__nand2_1 _39812_ (.A(_17438_),
    .B(_17439_),
    .Y(_17440_));
 sky130_fd_sc_hd__nor2_1 _39813_ (.A(_17433_),
    .B(_17251_),
    .Y(_17441_));
 sky130_fd_sc_hd__nand2_1 _39814_ (.A(_17440_),
    .B(_17441_),
    .Y(_17442_));
 sky130_fd_sc_hd__nand3b_4 _39815_ (.A_N(_17441_),
    .B(_17438_),
    .C(_17439_),
    .Y(_17443_));
 sky130_fd_sc_hd__nand2_4 _39816_ (.A(_17442_),
    .B(_17443_),
    .Y(_17444_));
 sky130_vsdinv _39817_ (.A(_17444_),
    .Y(_17445_));
 sky130_fd_sc_hd__o21ai_4 _39818_ (.A1(_17429_),
    .A2(_17430_),
    .B1(_17445_),
    .Y(_17446_));
 sky130_fd_sc_hd__a21oi_4 _39819_ (.A1(_17313_),
    .A2(_17315_),
    .B1(_17311_),
    .Y(_17447_));
 sky130_fd_sc_hd__nand2_1 _39820_ (.A(_17426_),
    .B(_17427_),
    .Y(_17448_));
 sky130_fd_sc_hd__and2_1 _39821_ (.A(_17306_),
    .B(_17281_),
    .X(_17449_));
 sky130_fd_sc_hd__nand2_4 _39822_ (.A(_17448_),
    .B(_17449_),
    .Y(_17450_));
 sky130_fd_sc_hd__nand3_4 _39823_ (.A(_17426_),
    .B(_17428_),
    .C(_17427_),
    .Y(_17451_));
 sky130_fd_sc_hd__nand3_4 _39824_ (.A(_17450_),
    .B(_17444_),
    .C(_17451_),
    .Y(_17452_));
 sky130_fd_sc_hd__nand3_4 _39825_ (.A(_17446_),
    .B(_17447_),
    .C(_17452_),
    .Y(_17453_));
 sky130_fd_sc_hd__o21ai_2 _39826_ (.A1(_17429_),
    .A2(_17430_),
    .B1(_17444_),
    .Y(_17454_));
 sky130_fd_sc_hd__nand3_2 _39827_ (.A(_17450_),
    .B(_17451_),
    .C(_17445_),
    .Y(_17455_));
 sky130_vsdinv _39828_ (.A(_17447_),
    .Y(_17456_));
 sky130_fd_sc_hd__nand3_4 _39829_ (.A(_17454_),
    .B(_17455_),
    .C(_17456_),
    .Y(_17457_));
 sky130_fd_sc_hd__o21ai_1 _39830_ (.A1(_17260_),
    .A2(_17261_),
    .B1(_17257_),
    .Y(_17458_));
 sky130_fd_sc_hd__or2_2 _39831_ (.A(_17237_),
    .B(_17458_),
    .X(_17459_));
 sky130_fd_sc_hd__nand2_2 _39832_ (.A(_17458_),
    .B(_17237_),
    .Y(_17460_));
 sky130_fd_sc_hd__clkbuf_2 _39833_ (.A(_17239_),
    .X(_17461_));
 sky130_fd_sc_hd__a21o_1 _39834_ (.A1(_17459_),
    .A2(_17460_),
    .B1(_17461_),
    .X(_17462_));
 sky130_fd_sc_hd__nand3_4 _39835_ (.A(_17459_),
    .B(_17239_),
    .C(_17460_),
    .Y(_17463_));
 sky130_fd_sc_hd__nand2_2 _39836_ (.A(_17462_),
    .B(_17463_),
    .Y(_17464_));
 sky130_fd_sc_hd__a21o_1 _39837_ (.A1(_17453_),
    .A2(_17457_),
    .B1(_17464_),
    .X(_17465_));
 sky130_fd_sc_hd__nand3_2 _39838_ (.A(_17453_),
    .B(_17457_),
    .C(_17464_),
    .Y(_17466_));
 sky130_fd_sc_hd__nand3b_4 _39839_ (.A_N(_17380_),
    .B(_17465_),
    .C(_17466_),
    .Y(_17467_));
 sky130_fd_sc_hd__and2_2 _39840_ (.A(_17462_),
    .B(_17463_),
    .X(_17468_));
 sky130_fd_sc_hd__a21o_1 _39841_ (.A1(_17453_),
    .A2(_17457_),
    .B1(_17468_),
    .X(_17469_));
 sky130_fd_sc_hd__nand3_4 _39842_ (.A(_17468_),
    .B(_17453_),
    .C(_17457_),
    .Y(_17470_));
 sky130_fd_sc_hd__nand3_4 _39843_ (.A(_17469_),
    .B(_17380_),
    .C(_17470_),
    .Y(_17471_));
 sky130_fd_sc_hd__nand2_1 _39844_ (.A(_17467_),
    .B(_17471_),
    .Y(_17472_));
 sky130_fd_sc_hd__nand2_1 _39845_ (.A(_17241_),
    .B(_17238_),
    .Y(_17473_));
 sky130_fd_sc_hd__or2_2 _39846_ (.A(_16835_),
    .B(_17473_),
    .X(_17474_));
 sky130_fd_sc_hd__nand2_2 _39847_ (.A(_17473_),
    .B(_17012_),
    .Y(_17475_));
 sky130_fd_sc_hd__buf_4 _39848_ (.A(_16841_),
    .X(_17476_));
 sky130_fd_sc_hd__a21oi_4 _39849_ (.A1(_17474_),
    .A2(_17475_),
    .B1(_17476_),
    .Y(_17477_));
 sky130_fd_sc_hd__and3_2 _39850_ (.A(_17474_),
    .B(_17476_),
    .C(_17475_),
    .X(_17478_));
 sky130_fd_sc_hd__nor2_8 _39851_ (.A(_17477_),
    .B(_17478_),
    .Y(_17479_));
 sky130_fd_sc_hd__nand2_4 _39852_ (.A(_17472_),
    .B(_17479_),
    .Y(_17480_));
 sky130_fd_sc_hd__nand3b_4 _39853_ (.A_N(_17479_),
    .B(_17467_),
    .C(_17471_),
    .Y(_17481_));
 sky130_vsdinv _39854_ (.A(_17329_),
    .Y(_17482_));
 sky130_fd_sc_hd__and2_1 _39855_ (.A(_17334_),
    .B(_17342_),
    .X(_17483_));
 sky130_fd_sc_hd__or2_4 _39856_ (.A(_17482_),
    .B(_17483_),
    .X(_17484_));
 sky130_fd_sc_hd__a21oi_4 _39857_ (.A1(_17480_),
    .A2(_17481_),
    .B1(_17484_),
    .Y(_17485_));
 sky130_fd_sc_hd__o211a_1 _39858_ (.A1(_17482_),
    .A2(_17483_),
    .B1(_17481_),
    .C1(_17480_),
    .X(_17486_));
 sky130_fd_sc_hd__nand2_1 _39859_ (.A(_17337_),
    .B(_17203_),
    .Y(_17487_));
 sky130_fd_sc_hd__nand2_2 _39860_ (.A(_17487_),
    .B(_17336_),
    .Y(_17488_));
 sky130_fd_sc_hd__nor2_8 _39861_ (.A(_16313_),
    .B(_17488_),
    .Y(_17489_));
 sky130_vsdinv _39862_ (.A(_17488_),
    .Y(_17490_));
 sky130_fd_sc_hd__nor2_8 _39863_ (.A(_16318_),
    .B(_17490_),
    .Y(_17491_));
 sky130_fd_sc_hd__nor2_8 _39864_ (.A(_17489_),
    .B(_17491_),
    .Y(_17492_));
 sky130_fd_sc_hd__o21ai_2 _39865_ (.A1(_17485_),
    .A2(_17486_),
    .B1(_17492_),
    .Y(_17493_));
 sky130_fd_sc_hd__a21o_1 _39866_ (.A1(_17480_),
    .A2(_17481_),
    .B1(_17484_),
    .X(_17494_));
 sky130_fd_sc_hd__nand3_4 _39867_ (.A(_17484_),
    .B(_17481_),
    .C(_17480_),
    .Y(_17495_));
 sky130_fd_sc_hd__nand3b_2 _39868_ (.A_N(_17492_),
    .B(_17494_),
    .C(_17495_),
    .Y(_17496_));
 sky130_fd_sc_hd__nand2_1 _39869_ (.A(_17349_),
    .B(_17359_),
    .Y(_17497_));
 sky130_fd_sc_hd__nand2_2 _39870_ (.A(_17497_),
    .B(_17344_),
    .Y(_17498_));
 sky130_fd_sc_hd__nand3_4 _39871_ (.A(_17493_),
    .B(_17496_),
    .C(_17498_),
    .Y(_17499_));
 sky130_fd_sc_hd__o22ai_4 _39872_ (.A1(_17489_),
    .A2(_17491_),
    .B1(_17485_),
    .B2(_17486_),
    .Y(_17500_));
 sky130_vsdinv _39873_ (.A(_17498_),
    .Y(_17501_));
 sky130_fd_sc_hd__nand3_2 _39874_ (.A(_17494_),
    .B(_17495_),
    .C(_17492_),
    .Y(_17502_));
 sky130_fd_sc_hd__nand3_4 _39875_ (.A(_17500_),
    .B(_17501_),
    .C(_17502_),
    .Y(_17503_));
 sky130_fd_sc_hd__a21oi_1 _39876_ (.A1(_17499_),
    .A2(_17503_),
    .B1(_17364_),
    .Y(_17504_));
 sky130_fd_sc_hd__and3_1 _39877_ (.A(_17499_),
    .B(_17503_),
    .C(_17364_),
    .X(_17505_));
 sky130_fd_sc_hd__o21ai_4 _39878_ (.A1(_17369_),
    .A2(_17370_),
    .B1(_17366_),
    .Y(_17506_));
 sky130_fd_sc_hd__o21bai_1 _39879_ (.A1(_17504_),
    .A2(_17505_),
    .B1_N(_17506_),
    .Y(_17507_));
 sky130_fd_sc_hd__nand2_2 _39880_ (.A(_17503_),
    .B(_17364_),
    .Y(_17508_));
 sky130_vsdinv _39881_ (.A(_17499_),
    .Y(_17509_));
 sky130_fd_sc_hd__a21o_1 _39882_ (.A1(_17499_),
    .A2(_17503_),
    .B1(_17364_),
    .X(_17510_));
 sky130_fd_sc_hd__o211ai_4 _39883_ (.A1(_17508_),
    .A2(_17509_),
    .B1(_17506_),
    .C1(_17510_),
    .Y(_17511_));
 sky130_fd_sc_hd__and2_1 _39884_ (.A(_17507_),
    .B(_17511_),
    .X(_17512_));
 sky130_fd_sc_hd__o2111a_1 _39885_ (.A1(_17368_),
    .A2(_17372_),
    .B1(_17228_),
    .C1(_17375_),
    .D1(_17223_),
    .X(_17513_));
 sky130_fd_sc_hd__nand2_1 _39886_ (.A(_17063_),
    .B(_17513_),
    .Y(_17514_));
 sky130_fd_sc_hd__o2111ai_4 _39887_ (.A1(_17368_),
    .A2(_17372_),
    .B1(_17228_),
    .C1(_17375_),
    .D1(_17223_),
    .Y(_17515_));
 sky130_fd_sc_hd__a2bb2oi_1 _39888_ (.A1_N(_17368_),
    .A2_N(_17372_),
    .B1(_17375_),
    .B2(_17378_),
    .Y(_17516_));
 sky130_fd_sc_hd__o21a_1 _39889_ (.A1(_17066_),
    .A2(_17515_),
    .B1(_17516_),
    .X(_17517_));
 sky130_fd_sc_hd__o21ai_4 _39890_ (.A1(_17514_),
    .A2(_16888_),
    .B1(_17517_),
    .Y(_17518_));
 sky130_fd_sc_hd__o2111ai_4 _39891_ (.A1(_17050_),
    .A2(_17062_),
    .B1(_16881_),
    .C1(_16878_),
    .D1(_17054_),
    .Y(_17519_));
 sky130_fd_sc_hd__nor2_2 _39892_ (.A(_17515_),
    .B(_17519_),
    .Y(_17520_));
 sky130_fd_sc_hd__nand2_1 _39893_ (.A(_17520_),
    .B(_16892_),
    .Y(_17521_));
 sky130_fd_sc_hd__a21oi_4 _39894_ (.A1(_16130_),
    .A2(_16134_),
    .B1(_17521_),
    .Y(_17522_));
 sky130_fd_sc_hd__nor2_2 _39895_ (.A(_17518_),
    .B(_17522_),
    .Y(_17523_));
 sky130_vsdinv _39896_ (.A(_17523_),
    .Y(_17524_));
 sky130_fd_sc_hd__or2_1 _39897_ (.A(_17512_),
    .B(_17524_),
    .X(_17525_));
 sky130_fd_sc_hd__nand2_1 _39898_ (.A(_17524_),
    .B(_17512_),
    .Y(_17526_));
 sky130_fd_sc_hd__and2_2 _39899_ (.A(_17525_),
    .B(_17526_),
    .X(_02675_));
 sky130_fd_sc_hd__o21ai_1 _39900_ (.A1(_17492_),
    .A2(_17485_),
    .B1(_17495_),
    .Y(_17527_));
 sky130_fd_sc_hd__a21oi_4 _39901_ (.A1(_17469_),
    .A2(_17470_),
    .B1(_17380_),
    .Y(_17528_));
 sky130_fd_sc_hd__o21ai_2 _39902_ (.A1(_17479_),
    .A2(_17528_),
    .B1(_17471_),
    .Y(_17529_));
 sky130_fd_sc_hd__a21boi_2 _39903_ (.A1(_17392_),
    .A2(_17404_),
    .B1_N(_17393_),
    .Y(_17530_));
 sky130_fd_sc_hd__o21a_2 _39904_ (.A1(_17382_),
    .A2(_17385_),
    .B1(_17383_),
    .X(_17531_));
 sky130_vsdinv _39905_ (.A(_17531_),
    .Y(_17532_));
 sky130_fd_sc_hd__nand2_2 _39906_ (.A(_19581_),
    .B(_19846_),
    .Y(_17533_));
 sky130_fd_sc_hd__or4_4 _39907_ (.A(_19852_),
    .B(_16352_),
    .C(_15817_),
    .D(_13260_),
    .X(_17534_));
 sky130_fd_sc_hd__a22o_1 _39908_ (.A1(_15821_),
    .A2(_15316_),
    .B1(_13855_),
    .B2(_11293_),
    .X(_17535_));
 sky130_fd_sc_hd__nand2_2 _39909_ (.A(_17534_),
    .B(_17535_),
    .Y(_17536_));
 sky130_fd_sc_hd__or2_2 _39910_ (.A(_17533_),
    .B(_17536_),
    .X(_17537_));
 sky130_fd_sc_hd__nand2_2 _39911_ (.A(_17536_),
    .B(_17533_),
    .Y(_17538_));
 sky130_fd_sc_hd__nand3_2 _39912_ (.A(_17532_),
    .B(_17537_),
    .C(_17538_),
    .Y(_17539_));
 sky130_fd_sc_hd__nand2_2 _39913_ (.A(_17537_),
    .B(_17538_),
    .Y(_17540_));
 sky130_fd_sc_hd__nand2_4 _39914_ (.A(_17540_),
    .B(_17531_),
    .Y(_17541_));
 sky130_fd_sc_hd__nand2_1 _39915_ (.A(_15806_),
    .B(_19831_),
    .Y(_17542_));
 sky130_fd_sc_hd__nand2_1 _39916_ (.A(_19589_),
    .B(_11582_),
    .Y(_17543_));
 sky130_fd_sc_hd__a32o_1 _39917_ (.A1(_15930_),
    .A2(_11582_),
    .A3(_11583_),
    .B1(_17395_),
    .B2(_17543_),
    .X(_17544_));
 sky130_fd_sc_hd__nor2_1 _39918_ (.A(_17542_),
    .B(_17544_),
    .Y(_17545_));
 sky130_fd_sc_hd__and2_1 _39919_ (.A(_17544_),
    .B(_17542_),
    .X(_17546_));
 sky130_fd_sc_hd__or2_2 _39920_ (.A(_17545_),
    .B(_17546_),
    .X(_17547_));
 sky130_fd_sc_hd__nand3_2 _39921_ (.A(_17539_),
    .B(_17541_),
    .C(_17547_),
    .Y(_17548_));
 sky130_fd_sc_hd__nand2_1 _39922_ (.A(_17540_),
    .B(_17532_),
    .Y(_17549_));
 sky130_fd_sc_hd__nand3_2 _39923_ (.A(_17537_),
    .B(_17531_),
    .C(_17538_),
    .Y(_17550_));
 sky130_vsdinv _39924_ (.A(_17547_),
    .Y(_17551_));
 sky130_fd_sc_hd__nand3_2 _39925_ (.A(_17549_),
    .B(_17550_),
    .C(_17551_),
    .Y(_17552_));
 sky130_fd_sc_hd__nand3_4 _39926_ (.A(_17530_),
    .B(_17548_),
    .C(_17552_),
    .Y(_17553_));
 sky130_fd_sc_hd__a21oi_1 _39927_ (.A1(_17386_),
    .A2(_17387_),
    .B1(_17390_),
    .Y(_17554_));
 sky130_fd_sc_hd__o21ai_2 _39928_ (.A1(_17400_),
    .A2(_17554_),
    .B1(_17393_),
    .Y(_17555_));
 sky130_fd_sc_hd__nand3_2 _39929_ (.A(_17539_),
    .B(_17541_),
    .C(_17551_),
    .Y(_17556_));
 sky130_fd_sc_hd__nand3_2 _39930_ (.A(_17549_),
    .B(_17550_),
    .C(_17547_),
    .Y(_17557_));
 sky130_fd_sc_hd__nand3_4 _39931_ (.A(_17555_),
    .B(_17556_),
    .C(_17557_),
    .Y(_17558_));
 sky130_fd_sc_hd__a31o_1 _39932_ (.A1(_19842_),
    .A2(_19846_),
    .A3(_16946_),
    .B1(_17398_),
    .X(_17559_));
 sky130_fd_sc_hd__nand2_2 _39933_ (.A(_11596_),
    .B(_14084_),
    .Y(_17560_));
 sky130_fd_sc_hd__or3_4 _39934_ (.A(_17560_),
    .B(_16940_),
    .C(_13007_),
    .X(_17561_));
 sky130_fd_sc_hd__o21ai_1 _39935_ (.A1(_16940_),
    .A2(_13007_),
    .B1(_17560_),
    .Y(_17562_));
 sky130_fd_sc_hd__nand2_1 _39936_ (.A(_17561_),
    .B(_17562_),
    .Y(_17563_));
 sky130_fd_sc_hd__nor2_2 _39937_ (.A(_17410_),
    .B(_17563_),
    .Y(_17564_));
 sky130_fd_sc_hd__nand2_1 _39938_ (.A(_17563_),
    .B(_17410_),
    .Y(_17565_));
 sky130_fd_sc_hd__and2b_1 _39939_ (.A_N(_17564_),
    .B(_17565_),
    .X(_17566_));
 sky130_fd_sc_hd__nor2_2 _39940_ (.A(_17559_),
    .B(_17566_),
    .Y(_17567_));
 sky130_vsdinv _39941_ (.A(_17567_),
    .Y(_17568_));
 sky130_fd_sc_hd__nand2_2 _39942_ (.A(_17414_),
    .B(_17411_),
    .Y(_17569_));
 sky130_vsdinv _39943_ (.A(_17569_),
    .Y(_17570_));
 sky130_fd_sc_hd__and3b_1 _39944_ (.A_N(_17564_),
    .B(_17559_),
    .C(_17565_),
    .X(_17571_));
 sky130_fd_sc_hd__inv_2 _39945_ (.A(_17571_),
    .Y(_17572_));
 sky130_fd_sc_hd__nand3_2 _39946_ (.A(_17568_),
    .B(_17570_),
    .C(_17572_),
    .Y(_17573_));
 sky130_fd_sc_hd__o21ai_2 _39947_ (.A1(_17571_),
    .A2(_17567_),
    .B1(_17569_),
    .Y(_17574_));
 sky130_fd_sc_hd__nand2_4 _39948_ (.A(_17573_),
    .B(_17574_),
    .Y(_17575_));
 sky130_fd_sc_hd__a21oi_2 _39949_ (.A1(_17553_),
    .A2(_17558_),
    .B1(_17575_),
    .Y(_17576_));
 sky130_fd_sc_hd__and3_1 _39950_ (.A(_17553_),
    .B(_17575_),
    .C(_17558_),
    .X(_17577_));
 sky130_fd_sc_hd__a21boi_2 _39951_ (.A1(_17425_),
    .A2(_17406_),
    .B1_N(_17409_),
    .Y(_17578_));
 sky130_fd_sc_hd__o21ai_4 _39952_ (.A1(_17576_),
    .A2(_17577_),
    .B1(_17578_),
    .Y(_17579_));
 sky130_fd_sc_hd__nand2_2 _39953_ (.A(_17427_),
    .B(_17409_),
    .Y(_17580_));
 sky130_fd_sc_hd__a21o_1 _39954_ (.A1(_17553_),
    .A2(_17558_),
    .B1(_17575_),
    .X(_17581_));
 sky130_fd_sc_hd__nand3_4 _39955_ (.A(_17553_),
    .B(_17575_),
    .C(_17558_),
    .Y(_17582_));
 sky130_fd_sc_hd__nand3_4 _39956_ (.A(_17580_),
    .B(_17581_),
    .C(_17582_),
    .Y(_17583_));
 sky130_fd_sc_hd__o21ai_1 _39957_ (.A1(_17422_),
    .A2(_17417_),
    .B1(_17423_),
    .Y(_17584_));
 sky130_fd_sc_hd__buf_4 _39958_ (.A(_17435_),
    .X(_17585_));
 sky130_fd_sc_hd__a21oi_4 _39959_ (.A1(_17434_),
    .A2(_17585_),
    .B1(_17436_),
    .Y(_17586_));
 sky130_fd_sc_hd__nand2_2 _39960_ (.A(_17584_),
    .B(_17586_),
    .Y(_17587_));
 sky130_fd_sc_hd__clkbuf_4 _39961_ (.A(_17437_),
    .X(_17588_));
 sky130_fd_sc_hd__o211ai_4 _39962_ (.A1(_17422_),
    .A2(_17417_),
    .B1(_17423_),
    .C1(_17588_),
    .Y(_17589_));
 sky130_fd_sc_hd__nand2_1 _39963_ (.A(_17587_),
    .B(_17589_),
    .Y(_17590_));
 sky130_vsdinv _39964_ (.A(_17585_),
    .Y(_17591_));
 sky130_fd_sc_hd__nand2_2 _39965_ (.A(_17590_),
    .B(_17591_),
    .Y(_17592_));
 sky130_fd_sc_hd__nand3_4 _39966_ (.A(_17587_),
    .B(_17589_),
    .C(_17585_),
    .Y(_17593_));
 sky130_fd_sc_hd__nand2_4 _39967_ (.A(_17592_),
    .B(_17593_),
    .Y(_17594_));
 sky130_fd_sc_hd__a21o_1 _39968_ (.A1(_17579_),
    .A2(_17583_),
    .B1(_17594_),
    .X(_17595_));
 sky130_fd_sc_hd__a21oi_4 _39969_ (.A1(_17450_),
    .A2(_17445_),
    .B1(_17430_),
    .Y(_17596_));
 sky130_fd_sc_hd__nand3_4 _39970_ (.A(_17579_),
    .B(_17583_),
    .C(_17594_),
    .Y(_17597_));
 sky130_fd_sc_hd__nand3_4 _39971_ (.A(_17595_),
    .B(_17596_),
    .C(_17597_),
    .Y(_17598_));
 sky130_vsdinv _39972_ (.A(_17592_),
    .Y(_17599_));
 sky130_vsdinv _39973_ (.A(_17593_),
    .Y(_17600_));
 sky130_fd_sc_hd__o2bb2ai_2 _39974_ (.A1_N(_17583_),
    .A2_N(_17579_),
    .B1(_17599_),
    .B2(_17600_),
    .Y(_17601_));
 sky130_fd_sc_hd__o21ai_2 _39975_ (.A1(_17444_),
    .A2(_17429_),
    .B1(_17451_),
    .Y(_17602_));
 sky130_fd_sc_hd__nand3b_4 _39976_ (.A_N(_17594_),
    .B(_17579_),
    .C(_17583_),
    .Y(_17603_));
 sky130_fd_sc_hd__nand3_4 _39977_ (.A(_17601_),
    .B(_17602_),
    .C(_17603_),
    .Y(_17604_));
 sky130_fd_sc_hd__nand2_2 _39978_ (.A(_17443_),
    .B(_17438_),
    .Y(_17605_));
 sky130_fd_sc_hd__nor2_4 _39979_ (.A(_17237_),
    .B(_17605_),
    .Y(_17606_));
 sky130_fd_sc_hd__buf_2 _39980_ (.A(_17237_),
    .X(_17607_));
 sky130_fd_sc_hd__nand2_1 _39981_ (.A(_17605_),
    .B(_17607_),
    .Y(_17608_));
 sky130_fd_sc_hd__nand2_2 _39982_ (.A(_17608_),
    .B(_17461_),
    .Y(_17609_));
 sky130_fd_sc_hd__a21o_1 _39983_ (.A1(_17166_),
    .A2(_17165_),
    .B1(_17605_),
    .X(_17610_));
 sky130_fd_sc_hd__nand2_1 _39984_ (.A(_17610_),
    .B(_17608_),
    .Y(_17611_));
 sky130_vsdinv _39985_ (.A(_17239_),
    .Y(_17612_));
 sky130_fd_sc_hd__buf_2 _39986_ (.A(_17612_),
    .X(_17613_));
 sky130_fd_sc_hd__nand2_2 _39987_ (.A(_17611_),
    .B(_17613_),
    .Y(_17614_));
 sky130_fd_sc_hd__o21ai_4 _39988_ (.A1(_17606_),
    .A2(_17609_),
    .B1(_17614_),
    .Y(_17615_));
 sky130_fd_sc_hd__a21o_1 _39989_ (.A1(_17598_),
    .A2(_17604_),
    .B1(_17615_),
    .X(_17616_));
 sky130_fd_sc_hd__a21oi_4 _39990_ (.A1(_17446_),
    .A2(_17452_),
    .B1(_17447_),
    .Y(_17617_));
 sky130_fd_sc_hd__a21oi_4 _39991_ (.A1(_17468_),
    .A2(_17453_),
    .B1(_17617_),
    .Y(_17618_));
 sky130_fd_sc_hd__nand3_4 _39992_ (.A(_17598_),
    .B(_17615_),
    .C(_17604_),
    .Y(_17619_));
 sky130_fd_sc_hd__nand3_4 _39993_ (.A(_17616_),
    .B(_17618_),
    .C(_17619_),
    .Y(_17620_));
 sky130_fd_sc_hd__a31oi_4 _39994_ (.A1(_17446_),
    .A2(_17447_),
    .A3(_17452_),
    .B1(_17464_),
    .Y(_17621_));
 sky130_fd_sc_hd__o21a_1 _39995_ (.A1(_17606_),
    .A2(_17609_),
    .B1(_17614_),
    .X(_17622_));
 sky130_fd_sc_hd__nand3_4 _39996_ (.A(_17622_),
    .B(_17598_),
    .C(_17604_),
    .Y(_17623_));
 sky130_fd_sc_hd__nor2_1 _39997_ (.A(_17606_),
    .B(_17609_),
    .Y(_17624_));
 sky130_vsdinv _39998_ (.A(_17614_),
    .Y(_17625_));
 sky130_fd_sc_hd__o2bb2ai_1 _39999_ (.A1_N(_17604_),
    .A2_N(_17598_),
    .B1(_17624_),
    .B2(_17625_),
    .Y(_17626_));
 sky130_fd_sc_hd__o211ai_4 _40000_ (.A1(_17617_),
    .A2(_17621_),
    .B1(_17623_),
    .C1(_17626_),
    .Y(_17627_));
 sky130_fd_sc_hd__a21o_1 _40001_ (.A1(_17463_),
    .A2(_17460_),
    .B1(_16478_),
    .X(_17628_));
 sky130_fd_sc_hd__nand3_2 _40002_ (.A(_17463_),
    .B(_16478_),
    .C(_17460_),
    .Y(_17629_));
 sky130_fd_sc_hd__nand2_4 _40003_ (.A(_17628_),
    .B(_17629_),
    .Y(_17630_));
 sky130_fd_sc_hd__xor2_4 _40004_ (.A(_17476_),
    .B(_17630_),
    .X(_17631_));
 sky130_fd_sc_hd__a21o_1 _40005_ (.A1(_17620_),
    .A2(_17627_),
    .B1(_17631_),
    .X(_17632_));
 sky130_fd_sc_hd__nand3_4 _40006_ (.A(_17631_),
    .B(_17620_),
    .C(_17627_),
    .Y(_17633_));
 sky130_fd_sc_hd__nand3_4 _40007_ (.A(_17529_),
    .B(_17632_),
    .C(_17633_),
    .Y(_17634_));
 sky130_fd_sc_hd__clkbuf_2 _40008_ (.A(_16484_),
    .X(_17635_));
 sky130_fd_sc_hd__nor2_1 _40009_ (.A(_17635_),
    .B(_17630_),
    .Y(_17636_));
 sky130_fd_sc_hd__and2_1 _40010_ (.A(_17630_),
    .B(_17635_),
    .X(_17637_));
 sky130_fd_sc_hd__nor2_1 _40011_ (.A(_17636_),
    .B(_17637_),
    .Y(_17638_));
 sky130_fd_sc_hd__nand3_2 _40012_ (.A(_17638_),
    .B(_17620_),
    .C(_17627_),
    .Y(_17639_));
 sky130_fd_sc_hd__o2bb2ai_1 _40013_ (.A1_N(_17627_),
    .A2_N(_17620_),
    .B1(_17637_),
    .B2(_17636_),
    .Y(_17640_));
 sky130_fd_sc_hd__o2111ai_4 _40014_ (.A1(_17479_),
    .A2(_17528_),
    .B1(_17471_),
    .C1(_17639_),
    .D1(_17640_),
    .Y(_17641_));
 sky130_fd_sc_hd__nand2_1 _40015_ (.A(_17474_),
    .B(_17635_),
    .Y(_17642_));
 sky130_fd_sc_hd__nand2_2 _40016_ (.A(_17642_),
    .B(_17475_),
    .Y(_17643_));
 sky130_fd_sc_hd__nor2_4 _40017_ (.A(_16313_),
    .B(_17643_),
    .Y(_17644_));
 sky130_vsdinv _40018_ (.A(_17643_),
    .Y(_17645_));
 sky130_fd_sc_hd__nor2_4 _40019_ (.A(_16318_),
    .B(_17645_),
    .Y(_17646_));
 sky130_fd_sc_hd__nor2_4 _40020_ (.A(_17644_),
    .B(_17646_),
    .Y(_17647_));
 sky130_fd_sc_hd__a21bo_1 _40021_ (.A1(_17634_),
    .A2(_17641_),
    .B1_N(_17647_),
    .X(_17648_));
 sky130_fd_sc_hd__nand3b_1 _40022_ (.A_N(_17647_),
    .B(_17634_),
    .C(_17641_),
    .Y(_17649_));
 sky130_fd_sc_hd__nand3_2 _40023_ (.A(_17527_),
    .B(_17648_),
    .C(_17649_),
    .Y(_17650_));
 sky130_fd_sc_hd__nand3_2 _40024_ (.A(_17634_),
    .B(_17641_),
    .C(_17647_),
    .Y(_17651_));
 sky130_fd_sc_hd__o2bb2ai_2 _40025_ (.A1_N(_17641_),
    .A2_N(_17634_),
    .B1(_17644_),
    .B2(_17646_),
    .Y(_17652_));
 sky130_fd_sc_hd__o2111ai_4 _40026_ (.A1(_17492_),
    .A2(_17485_),
    .B1(_17495_),
    .C1(_17651_),
    .D1(_17652_),
    .Y(_17653_));
 sky130_fd_sc_hd__nor2_1 _40027_ (.A(_16515_),
    .B(_17490_),
    .Y(_17654_));
 sky130_fd_sc_hd__a21oi_1 _40028_ (.A1(_17650_),
    .A2(_17653_),
    .B1(_17654_),
    .Y(_17655_));
 sky130_fd_sc_hd__and3_1 _40029_ (.A(_17650_),
    .B(_17653_),
    .C(_17654_),
    .X(_17656_));
 sky130_fd_sc_hd__a211o_1 _40030_ (.A1(_17499_),
    .A2(_17508_),
    .B1(_17655_),
    .C1(_17656_),
    .X(_17657_));
 sky130_fd_sc_hd__a21oi_1 _40031_ (.A1(_17364_),
    .A2(_17503_),
    .B1(_17509_),
    .Y(_17658_));
 sky130_fd_sc_hd__o21ai_1 _40032_ (.A1(_17655_),
    .A2(_17656_),
    .B1(_17658_),
    .Y(_17659_));
 sky130_fd_sc_hd__and2_2 _40033_ (.A(_17657_),
    .B(_17659_),
    .X(_17660_));
 sky130_fd_sc_hd__nand2_2 _40034_ (.A(_17526_),
    .B(_17511_),
    .Y(_17661_));
 sky130_fd_sc_hd__xor2_4 _40035_ (.A(_17660_),
    .B(_17661_),
    .X(_02676_));
 sky130_fd_sc_hd__nor2_2 _40036_ (.A(net410),
    .B(_17645_),
    .Y(_17662_));
 sky130_vsdinv _40037_ (.A(_17662_),
    .Y(_17663_));
 sky130_fd_sc_hd__nand2_1 _40038_ (.A(_17593_),
    .B(_17587_),
    .Y(_17664_));
 sky130_fd_sc_hd__or2_2 _40039_ (.A(_17607_),
    .B(_17664_),
    .X(_17665_));
 sky130_fd_sc_hd__nand2_1 _40040_ (.A(_17664_),
    .B(_17607_),
    .Y(_17666_));
 sky130_fd_sc_hd__nand3_1 _40041_ (.A(_17665_),
    .B(_17461_),
    .C(_17666_),
    .Y(_17667_));
 sky130_vsdinv _40042_ (.A(_17667_),
    .Y(_17668_));
 sky130_fd_sc_hd__nand2_1 _40043_ (.A(_17665_),
    .B(_17666_),
    .Y(_17669_));
 sky130_fd_sc_hd__nand2_1 _40044_ (.A(_17669_),
    .B(_17613_),
    .Y(_17670_));
 sky130_vsdinv _40045_ (.A(_17670_),
    .Y(_17671_));
 sky130_fd_sc_hd__nand3_2 _40046_ (.A(_17568_),
    .B(_17569_),
    .C(_17572_),
    .Y(_17672_));
 sky130_fd_sc_hd__a21o_1 _40047_ (.A1(_17672_),
    .A2(_17572_),
    .B1(_17588_),
    .X(_17673_));
 sky130_fd_sc_hd__nand3_2 _40048_ (.A(_17672_),
    .B(_17588_),
    .C(_17572_),
    .Y(_17674_));
 sky130_fd_sc_hd__nand3_4 _40049_ (.A(_17673_),
    .B(_17585_),
    .C(_17674_),
    .Y(_17675_));
 sky130_vsdinv _40050_ (.A(_17675_),
    .Y(_17676_));
 sky130_fd_sc_hd__o211a_1 _40051_ (.A1(_17567_),
    .A2(_17570_),
    .B1(_17572_),
    .C1(_17588_),
    .X(_17677_));
 sky130_fd_sc_hd__a21oi_1 _40052_ (.A1(_17672_),
    .A2(_17572_),
    .B1(_17588_),
    .Y(_17678_));
 sky130_fd_sc_hd__o21ai_2 _40053_ (.A1(_17677_),
    .A2(_17678_),
    .B1(_17591_),
    .Y(_17679_));
 sky130_vsdinv _40054_ (.A(_17679_),
    .Y(_17680_));
 sky130_fd_sc_hd__nor2_2 _40055_ (.A(_17531_),
    .B(_17540_),
    .Y(_17681_));
 sky130_fd_sc_hd__a21oi_4 _40056_ (.A1(_17541_),
    .A2(_17551_),
    .B1(_17681_),
    .Y(_17682_));
 sky130_fd_sc_hd__nand2_1 _40057_ (.A(_19594_),
    .B(_19828_),
    .Y(_17683_));
 sky130_fd_sc_hd__o22a_1 _40058_ (.A1(_16159_),
    .A2(_11206_),
    .B1(_15834_),
    .B2(_13309_),
    .X(_17684_));
 sky130_fd_sc_hd__a31o_1 _40059_ (.A1(_19832_),
    .A2(_19836_),
    .A3(_16946_),
    .B1(_17684_),
    .X(_17685_));
 sky130_fd_sc_hd__nor2_4 _40060_ (.A(_17683_),
    .B(_17685_),
    .Y(_17686_));
 sky130_fd_sc_hd__and2_2 _40061_ (.A(_17685_),
    .B(_17683_),
    .X(_17687_));
 sky130_fd_sc_hd__nor2_8 _40062_ (.A(_17686_),
    .B(_17687_),
    .Y(_17688_));
 sky130_fd_sc_hd__o21ai_2 _40063_ (.A1(_17533_),
    .A2(_17536_),
    .B1(_17534_),
    .Y(_17689_));
 sky130_fd_sc_hd__nand2_1 _40064_ (.A(_19580_),
    .B(_19842_),
    .Y(_17690_));
 sky130_vsdinv _40065_ (.A(_17690_),
    .Y(_17691_));
 sky130_fd_sc_hd__or4_4 _40066_ (.A(_15316_),
    .B(_18476_),
    .C(_16353_),
    .D(_13900_),
    .X(_17692_));
 sky130_fd_sc_hd__a22o_1 _40067_ (.A1(_19578_),
    .A2(_19845_),
    .B1(_13260_),
    .B2(_11293_),
    .X(_17693_));
 sky130_fd_sc_hd__nand2_2 _40068_ (.A(_17692_),
    .B(_17693_),
    .Y(_17694_));
 sky130_fd_sc_hd__or2_1 _40069_ (.A(_17691_),
    .B(_17694_),
    .X(_17695_));
 sky130_fd_sc_hd__nand2_1 _40070_ (.A(_17694_),
    .B(_17691_),
    .Y(_17696_));
 sky130_fd_sc_hd__nand3b_4 _40071_ (.A_N(_17689_),
    .B(_17695_),
    .C(_17696_),
    .Y(_17697_));
 sky130_fd_sc_hd__or2_1 _40072_ (.A(_17690_),
    .B(_17694_),
    .X(_17698_));
 sky130_fd_sc_hd__nand2_1 _40073_ (.A(_17694_),
    .B(_17690_),
    .Y(_17699_));
 sky130_fd_sc_hd__nand3_4 _40074_ (.A(_17698_),
    .B(_17689_),
    .C(_17699_),
    .Y(_17700_));
 sky130_fd_sc_hd__nand3b_4 _40075_ (.A_N(_17688_),
    .B(_17697_),
    .C(_17700_),
    .Y(_17701_));
 sky130_fd_sc_hd__a21bo_1 _40076_ (.A1(_17697_),
    .A2(_17700_),
    .B1_N(_17688_),
    .X(_17702_));
 sky130_fd_sc_hd__nand3_4 _40077_ (.A(_17682_),
    .B(_17701_),
    .C(_17702_),
    .Y(_17703_));
 sky130_fd_sc_hd__a21o_1 _40078_ (.A1(_17541_),
    .A2(_17551_),
    .B1(_17681_),
    .X(_17704_));
 sky130_fd_sc_hd__nand3_4 _40079_ (.A(_17697_),
    .B(_17700_),
    .C(_17688_),
    .Y(_17705_));
 sky130_fd_sc_hd__a21o_1 _40080_ (.A1(_17697_),
    .A2(_17700_),
    .B1(_17688_),
    .X(_17706_));
 sky130_fd_sc_hd__nand3_4 _40081_ (.A(_17704_),
    .B(_17705_),
    .C(_17706_),
    .Y(_17707_));
 sky130_vsdinv _40082_ (.A(_17561_),
    .Y(_17708_));
 sky130_fd_sc_hd__nor2_4 _40083_ (.A(_17708_),
    .B(_17564_),
    .Y(_17709_));
 sky130_fd_sc_hd__a31o_1 _40084_ (.A1(_19837_),
    .A2(_19842_),
    .A3(_16946_),
    .B1(_17545_),
    .X(_17710_));
 sky130_fd_sc_hd__nand2_2 _40085_ (.A(_12614_),
    .B(_13514_),
    .Y(_17711_));
 sky130_fd_sc_hd__or2_2 _40086_ (.A(_17711_),
    .B(_15957_),
    .X(_17712_));
 sky130_fd_sc_hd__nand2_1 _40087_ (.A(_17560_),
    .B(_17711_),
    .Y(_17713_));
 sky130_fd_sc_hd__nand2_1 _40088_ (.A(_17712_),
    .B(_17713_),
    .Y(_17714_));
 sky130_fd_sc_hd__or2_1 _40089_ (.A(_17410_),
    .B(_17714_),
    .X(_17715_));
 sky130_fd_sc_hd__nand2_1 _40090_ (.A(_17714_),
    .B(_17410_),
    .Y(_17716_));
 sky130_fd_sc_hd__and2_2 _40091_ (.A(_17715_),
    .B(_17716_),
    .X(_17717_));
 sky130_fd_sc_hd__or2_4 _40092_ (.A(_17710_),
    .B(_17717_),
    .X(_17718_));
 sky130_fd_sc_hd__nand2_4 _40093_ (.A(_17717_),
    .B(_17710_),
    .Y(_17719_));
 sky130_fd_sc_hd__nand2_2 _40094_ (.A(_17718_),
    .B(_17719_),
    .Y(_17720_));
 sky130_fd_sc_hd__nor2_4 _40095_ (.A(_17709_),
    .B(_17720_),
    .Y(_17721_));
 sky130_fd_sc_hd__a21boi_4 _40096_ (.A1(_17718_),
    .A2(_17719_),
    .B1_N(_17709_),
    .Y(_17722_));
 sky130_fd_sc_hd__o2bb2ai_2 _40097_ (.A1_N(_17703_),
    .A2_N(_17707_),
    .B1(_17721_),
    .B2(_17722_),
    .Y(_17723_));
 sky130_fd_sc_hd__a21o_1 _40098_ (.A1(_17718_),
    .A2(_17719_),
    .B1(_17709_),
    .X(_17724_));
 sky130_fd_sc_hd__nand3_1 _40099_ (.A(_17718_),
    .B(_17709_),
    .C(_17719_),
    .Y(_17725_));
 sky130_fd_sc_hd__nand2_2 _40100_ (.A(_17724_),
    .B(_17725_),
    .Y(_17726_));
 sky130_fd_sc_hd__nand3_2 _40101_ (.A(_17707_),
    .B(_17726_),
    .C(_17703_),
    .Y(_17727_));
 sky130_fd_sc_hd__nand2_2 _40102_ (.A(_17582_),
    .B(_17558_),
    .Y(_17728_));
 sky130_fd_sc_hd__a21oi_4 _40103_ (.A1(_17723_),
    .A2(_17727_),
    .B1(_17728_),
    .Y(_17729_));
 sky130_fd_sc_hd__a21boi_4 _40104_ (.A1(_17553_),
    .A2(_17575_),
    .B1_N(_17558_),
    .Y(_17730_));
 sky130_fd_sc_hd__a2bb2oi_4 _40105_ (.A1_N(_17721_),
    .A2_N(_17722_),
    .B1(_17703_),
    .B2(_17707_),
    .Y(_17731_));
 sky130_fd_sc_hd__and3_4 _40106_ (.A(_17707_),
    .B(_17726_),
    .C(_17703_),
    .X(_17732_));
 sky130_fd_sc_hd__nor3_4 _40107_ (.A(_17730_),
    .B(_17731_),
    .C(_17732_),
    .Y(_17733_));
 sky130_fd_sc_hd__o22ai_4 _40108_ (.A1(_17676_),
    .A2(_17680_),
    .B1(_17729_),
    .B2(_17733_),
    .Y(_17734_));
 sky130_fd_sc_hd__nand2_2 _40109_ (.A(_17723_),
    .B(_17728_),
    .Y(_17735_));
 sky130_fd_sc_hd__and2_1 _40110_ (.A(_17679_),
    .B(_17675_),
    .X(_17736_));
 sky130_fd_sc_hd__o21ai_2 _40111_ (.A1(_17731_),
    .A2(_17732_),
    .B1(_17730_),
    .Y(_17737_));
 sky130_fd_sc_hd__o211ai_4 _40112_ (.A1(_17732_),
    .A2(_17735_),
    .B1(_17736_),
    .C1(_17737_),
    .Y(_17738_));
 sky130_fd_sc_hd__a21oi_2 _40113_ (.A1(_17581_),
    .A2(_17582_),
    .B1(_17580_),
    .Y(_17739_));
 sky130_fd_sc_hd__o21ai_4 _40114_ (.A1(_17594_),
    .A2(_17739_),
    .B1(_17583_),
    .Y(_17740_));
 sky130_fd_sc_hd__a21oi_4 _40115_ (.A1(_17734_),
    .A2(_17738_),
    .B1(_17740_),
    .Y(_17741_));
 sky130_fd_sc_hd__and3_1 _40116_ (.A(_17734_),
    .B(_17738_),
    .C(_17740_),
    .X(_17742_));
 sky130_fd_sc_hd__o22ai_4 _40117_ (.A1(_17668_),
    .A2(_17671_),
    .B1(_17741_),
    .B2(_17742_),
    .Y(_17743_));
 sky130_fd_sc_hd__nand2_1 _40118_ (.A(_17670_),
    .B(_17667_),
    .Y(_17744_));
 sky130_fd_sc_hd__a21o_1 _40119_ (.A1(_17734_),
    .A2(_17738_),
    .B1(_17740_),
    .X(_17745_));
 sky130_fd_sc_hd__nand3_4 _40120_ (.A(_17734_),
    .B(_17738_),
    .C(_17740_),
    .Y(_17746_));
 sky130_fd_sc_hd__nand3b_4 _40121_ (.A_N(_17744_),
    .B(_17745_),
    .C(_17746_),
    .Y(_17747_));
 sky130_fd_sc_hd__and3_1 _40122_ (.A(_17601_),
    .B(_17602_),
    .C(_17603_),
    .X(_17748_));
 sky130_fd_sc_hd__a21o_2 _40123_ (.A1(_17598_),
    .A2(_17622_),
    .B1(_17748_),
    .X(_17749_));
 sky130_fd_sc_hd__a21oi_4 _40124_ (.A1(_17743_),
    .A2(_17747_),
    .B1(_17749_),
    .Y(_17750_));
 sky130_fd_sc_hd__a31oi_1 _40125_ (.A1(_17596_),
    .A2(_17597_),
    .A3(_17595_),
    .B1(_17615_),
    .Y(_17751_));
 sky130_fd_sc_hd__o211a_1 _40126_ (.A1(_17748_),
    .A2(_17751_),
    .B1(_17747_),
    .C1(_17743_),
    .X(_17752_));
 sky130_vsdinv _40127_ (.A(_17608_),
    .Y(_17753_));
 sky130_fd_sc_hd__nor2_1 _40128_ (.A(_17612_),
    .B(_17606_),
    .Y(_17754_));
 sky130_fd_sc_hd__or3_4 _40129_ (.A(_16835_),
    .B(_17753_),
    .C(_17754_),
    .X(_17755_));
 sky130_fd_sc_hd__o21ai_2 _40130_ (.A1(_17753_),
    .A2(_17754_),
    .B1(_17012_),
    .Y(_17756_));
 sky130_fd_sc_hd__a21o_1 _40131_ (.A1(_17755_),
    .A2(_17756_),
    .B1(_17203_),
    .X(_17757_));
 sky130_fd_sc_hd__nand3_2 _40132_ (.A(_17755_),
    .B(_17756_),
    .C(_17203_),
    .Y(_17758_));
 sky130_fd_sc_hd__nand2_2 _40133_ (.A(_17757_),
    .B(_17758_),
    .Y(_17759_));
 sky130_fd_sc_hd__o21ai_4 _40134_ (.A1(_17750_),
    .A2(_17752_),
    .B1(_17759_),
    .Y(_17760_));
 sky130_fd_sc_hd__a21o_1 _40135_ (.A1(_17743_),
    .A2(_17747_),
    .B1(_17749_),
    .X(_17761_));
 sky130_fd_sc_hd__and2_1 _40136_ (.A(_17757_),
    .B(_17758_),
    .X(_17762_));
 sky130_fd_sc_hd__nand3_4 _40137_ (.A(_17749_),
    .B(_17743_),
    .C(_17747_),
    .Y(_17763_));
 sky130_fd_sc_hd__nand3_4 _40138_ (.A(_17761_),
    .B(_17762_),
    .C(_17763_),
    .Y(_17764_));
 sky130_fd_sc_hd__a21oi_1 _40139_ (.A1(_17616_),
    .A2(_17619_),
    .B1(_17618_),
    .Y(_17765_));
 sky130_fd_sc_hd__a21o_2 _40140_ (.A1(_17631_),
    .A2(_17620_),
    .B1(_17765_),
    .X(_17766_));
 sky130_fd_sc_hd__a21oi_4 _40141_ (.A1(_17760_),
    .A2(_17764_),
    .B1(_17766_),
    .Y(_17767_));
 sky130_fd_sc_hd__and3_1 _40142_ (.A(_17760_),
    .B(_17766_),
    .C(_17764_),
    .X(_17768_));
 sky130_fd_sc_hd__o21a_2 _40143_ (.A1(_17476_),
    .A2(_17630_),
    .B1(_17628_),
    .X(_17769_));
 sky130_fd_sc_hd__or2_1 _40144_ (.A(_16675_),
    .B(_17769_),
    .X(_17770_));
 sky130_fd_sc_hd__nand2_1 _40145_ (.A(_17769_),
    .B(_16318_),
    .Y(_17771_));
 sky130_fd_sc_hd__nand2_2 _40146_ (.A(_17770_),
    .B(_17771_),
    .Y(_17772_));
 sky130_vsdinv _40147_ (.A(_17772_),
    .Y(_17773_));
 sky130_fd_sc_hd__o21ai_2 _40148_ (.A1(_17767_),
    .A2(_17768_),
    .B1(_17773_),
    .Y(_17774_));
 sky130_fd_sc_hd__nand2_1 _40149_ (.A(_17760_),
    .B(_17764_),
    .Y(_17775_));
 sky130_vsdinv _40150_ (.A(_17766_),
    .Y(_17776_));
 sky130_fd_sc_hd__nand2_2 _40151_ (.A(_17775_),
    .B(_17776_),
    .Y(_17777_));
 sky130_fd_sc_hd__nand3_4 _40152_ (.A(_17760_),
    .B(_17764_),
    .C(_17766_),
    .Y(_17778_));
 sky130_fd_sc_hd__nand3_4 _40153_ (.A(_17777_),
    .B(_17778_),
    .C(_17772_),
    .Y(_17779_));
 sky130_fd_sc_hd__a21oi_2 _40154_ (.A1(_17632_),
    .A2(_17633_),
    .B1(_17529_),
    .Y(_17780_));
 sky130_fd_sc_hd__o21ai_2 _40155_ (.A1(_17647_),
    .A2(_17780_),
    .B1(_17634_),
    .Y(_17781_));
 sky130_fd_sc_hd__nand3_4 _40156_ (.A(_17774_),
    .B(_17779_),
    .C(_17781_),
    .Y(_17782_));
 sky130_fd_sc_hd__o21ai_2 _40157_ (.A1(_17767_),
    .A2(_17768_),
    .B1(_17772_),
    .Y(_17783_));
 sky130_fd_sc_hd__o21a_1 _40158_ (.A1(_17647_),
    .A2(_17780_),
    .B1(_17634_),
    .X(_17784_));
 sky130_fd_sc_hd__nand3_4 _40159_ (.A(_17777_),
    .B(_17778_),
    .C(_17773_),
    .Y(_17785_));
 sky130_fd_sc_hd__nand3_4 _40160_ (.A(_17783_),
    .B(_17784_),
    .C(_17785_),
    .Y(_17786_));
 sky130_fd_sc_hd__nand2_2 _40161_ (.A(_17782_),
    .B(_17786_),
    .Y(_17787_));
 sky130_fd_sc_hd__nor2_4 _40162_ (.A(_17663_),
    .B(_17787_),
    .Y(_17788_));
 sky130_fd_sc_hd__clkbuf_4 _40163_ (.A(_16515_),
    .X(_17789_));
 sky130_fd_sc_hd__o2bb2ai_1 _40164_ (.A1_N(_17782_),
    .A2_N(_17786_),
    .B1(_17789_),
    .B2(_17645_),
    .Y(_17790_));
 sky130_fd_sc_hd__nand2_1 _40165_ (.A(_17653_),
    .B(_17654_),
    .Y(_17791_));
 sky130_fd_sc_hd__nand2_1 _40166_ (.A(_17791_),
    .B(_17650_),
    .Y(_17792_));
 sky130_fd_sc_hd__nand2_2 _40167_ (.A(_17790_),
    .B(_17792_),
    .Y(_17793_));
 sky130_fd_sc_hd__nand2_1 _40168_ (.A(_17787_),
    .B(_17662_),
    .Y(_17794_));
 sky130_fd_sc_hd__nand3_1 _40169_ (.A(_17782_),
    .B(_17786_),
    .C(_17663_),
    .Y(_17795_));
 sky130_fd_sc_hd__nand3b_2 _40170_ (.A_N(_17792_),
    .B(_17794_),
    .C(_17795_),
    .Y(_17796_));
 sky130_fd_sc_hd__o21a_2 _40171_ (.A1(_17788_),
    .A2(_17793_),
    .B1(_17796_),
    .X(_17797_));
 sky130_fd_sc_hd__nand2_1 _40172_ (.A(_17508_),
    .B(_17499_),
    .Y(_17798_));
 sky130_fd_sc_hd__o2bb2ai_1 _40173_ (.A1_N(_17650_),
    .A2_N(_17653_),
    .B1(_17789_),
    .B2(_17490_),
    .Y(_17799_));
 sky130_fd_sc_hd__nand2_1 _40174_ (.A(_17798_),
    .B(_17799_),
    .Y(_17800_));
 sky130_fd_sc_hd__o2111a_1 _40175_ (.A1(_17656_),
    .A2(_17800_),
    .B1(_17511_),
    .C1(_17659_),
    .D1(_17507_),
    .X(_17801_));
 sky130_vsdinv _40176_ (.A(_17801_),
    .Y(_17802_));
 sky130_vsdinv _40177_ (.A(_17659_),
    .Y(_17803_));
 sky130_fd_sc_hd__a21oi_4 _40178_ (.A1(_17657_),
    .A2(_17511_),
    .B1(_17803_),
    .Y(_17804_));
 sky130_fd_sc_hd__o21bai_4 _40179_ (.A1(_17802_),
    .A2(_17523_),
    .B1_N(_17804_),
    .Y(_17805_));
 sky130_fd_sc_hd__xor2_4 _40180_ (.A(_17797_),
    .B(_17805_),
    .X(_02677_));
 sky130_fd_sc_hd__buf_2 _40181_ (.A(_17635_),
    .X(_17806_));
 sky130_fd_sc_hd__a21boi_4 _40182_ (.A1(_17755_),
    .A2(_17806_),
    .B1_N(_17756_),
    .Y(_17807_));
 sky130_fd_sc_hd__nor2_8 _40183_ (.A(_14331_),
    .B(_17807_),
    .Y(_17808_));
 sky130_fd_sc_hd__and3_1 _40184_ (.A(_17758_),
    .B(_16313_),
    .C(_17756_),
    .X(_17809_));
 sky130_fd_sc_hd__o21a_1 _40185_ (.A1(_17690_),
    .A2(_17694_),
    .B1(_17692_),
    .X(_17810_));
 sky130_vsdinv _40186_ (.A(_17810_),
    .Y(_17811_));
 sky130_fd_sc_hd__nor2_1 _40187_ (.A(_15814_),
    .B(_15780_),
    .Y(_17812_));
 sky130_vsdinv _40188_ (.A(_17812_),
    .Y(_17813_));
 sky130_fd_sc_hd__or4_4 _40189_ (.A(_13248_),
    .B(_16352_),
    .C(_15817_),
    .D(_12902_),
    .X(_17814_));
 sky130_fd_sc_hd__a22o_1 _40190_ (.A1(_15821_),
    .A2(_11583_),
    .B1(_13900_),
    .B2(_11293_),
    .X(_17815_));
 sky130_fd_sc_hd__nand2_1 _40191_ (.A(_17814_),
    .B(_17815_),
    .Y(_17816_));
 sky130_fd_sc_hd__or2_1 _40192_ (.A(_17813_),
    .B(_17816_),
    .X(_17817_));
 sky130_fd_sc_hd__buf_2 _40193_ (.A(_17817_),
    .X(_17818_));
 sky130_fd_sc_hd__nand2_2 _40194_ (.A(_17816_),
    .B(_17813_),
    .Y(_17819_));
 sky130_fd_sc_hd__nand3_4 _40195_ (.A(_17811_),
    .B(_17818_),
    .C(_17819_),
    .Y(_17820_));
 sky130_fd_sc_hd__nand2_1 _40196_ (.A(_17818_),
    .B(_17819_),
    .Y(_17821_));
 sky130_fd_sc_hd__nand2_2 _40197_ (.A(_17821_),
    .B(_17810_),
    .Y(_17822_));
 sky130_fd_sc_hd__nand2_1 _40198_ (.A(_14218_),
    .B(_19594_),
    .Y(_17823_));
 sky130_vsdinv _40199_ (.A(_17823_),
    .Y(_17824_));
 sky130_fd_sc_hd__and4_1 _40200_ (.A(_19585_),
    .B(_19589_),
    .C(_19827_),
    .D(_19831_),
    .X(_17825_));
 sky130_fd_sc_hd__o22a_1 _40201_ (.A1(_16159_),
    .A2(_17288_),
    .B1(_15834_),
    .B2(_17245_),
    .X(_17826_));
 sky130_fd_sc_hd__nor2_1 _40202_ (.A(_17825_),
    .B(_17826_),
    .Y(_17827_));
 sky130_fd_sc_hd__or2_1 _40203_ (.A(_17824_),
    .B(_17827_),
    .X(_17828_));
 sky130_fd_sc_hd__buf_2 _40204_ (.A(_17824_),
    .X(_17829_));
 sky130_fd_sc_hd__nand2_1 _40205_ (.A(_17827_),
    .B(_17829_),
    .Y(_17830_));
 sky130_fd_sc_hd__nand2_2 _40206_ (.A(_17828_),
    .B(_17830_),
    .Y(_17831_));
 sky130_fd_sc_hd__nand3_2 _40207_ (.A(_17820_),
    .B(_17822_),
    .C(_17831_),
    .Y(_17832_));
 sky130_fd_sc_hd__a21o_1 _40208_ (.A1(_17818_),
    .A2(_17819_),
    .B1(_17810_),
    .X(_17833_));
 sky130_fd_sc_hd__nand3_2 _40209_ (.A(_17818_),
    .B(_17810_),
    .C(_17819_),
    .Y(_17834_));
 sky130_vsdinv _40210_ (.A(_17831_),
    .Y(_17835_));
 sky130_fd_sc_hd__nand3_2 _40211_ (.A(_17833_),
    .B(_17834_),
    .C(_17835_),
    .Y(_17836_));
 sky130_fd_sc_hd__a21boi_2 _40212_ (.A1(_17697_),
    .A2(_17688_),
    .B1_N(_17700_),
    .Y(_17837_));
 sky130_fd_sc_hd__nand3_4 _40213_ (.A(_17832_),
    .B(_17836_),
    .C(_17837_),
    .Y(_17838_));
 sky130_fd_sc_hd__nand2_1 _40214_ (.A(_17705_),
    .B(_17700_),
    .Y(_17839_));
 sky130_fd_sc_hd__nand3_4 _40215_ (.A(_17820_),
    .B(_17822_),
    .C(_17835_),
    .Y(_17840_));
 sky130_fd_sc_hd__nand3_2 _40216_ (.A(_17833_),
    .B(_17834_),
    .C(_17831_),
    .Y(_17841_));
 sky130_fd_sc_hd__nand3_4 _40217_ (.A(_17839_),
    .B(_17840_),
    .C(_17841_),
    .Y(_17842_));
 sky130_vsdinv _40218_ (.A(_17712_),
    .Y(_17843_));
 sky130_vsdinv _40219_ (.A(_17715_),
    .Y(_17844_));
 sky130_fd_sc_hd__nor2_4 _40220_ (.A(_17843_),
    .B(_17844_),
    .Y(_17845_));
 sky130_fd_sc_hd__clkbuf_2 _40221_ (.A(_17845_),
    .X(_17846_));
 sky130_fd_sc_hd__a31o_1 _40222_ (.A1(_19832_),
    .A2(_19837_),
    .A3(_16946_),
    .B1(_17686_),
    .X(_17847_));
 sky130_fd_sc_hd__a21o_1 _40223_ (.A1(_17715_),
    .A2(_17716_),
    .B1(_17847_),
    .X(_17848_));
 sky130_fd_sc_hd__nand2_2 _40224_ (.A(_17847_),
    .B(_17717_),
    .Y(_17849_));
 sky130_fd_sc_hd__nand2_2 _40225_ (.A(_17848_),
    .B(_17849_),
    .Y(_17850_));
 sky130_fd_sc_hd__nor2_1 _40226_ (.A(_17846_),
    .B(_17850_),
    .Y(_17851_));
 sky130_fd_sc_hd__and2_1 _40227_ (.A(_17850_),
    .B(_17845_),
    .X(_17852_));
 sky130_fd_sc_hd__o2bb2ai_2 _40228_ (.A1_N(_17838_),
    .A2_N(_17842_),
    .B1(_17851_),
    .B2(_17852_),
    .Y(_17853_));
 sky130_fd_sc_hd__a21oi_2 _40229_ (.A1(_17848_),
    .A2(_17849_),
    .B1(_17846_),
    .Y(_17854_));
 sky130_vsdinv _40230_ (.A(_17845_),
    .Y(_17855_));
 sky130_fd_sc_hd__nor2_2 _40231_ (.A(_17855_),
    .B(_17850_),
    .Y(_17856_));
 sky130_fd_sc_hd__o211ai_4 _40232_ (.A1(_17854_),
    .A2(_17856_),
    .B1(_17838_),
    .C1(_17842_),
    .Y(_17857_));
 sky130_fd_sc_hd__nand2_1 _40233_ (.A(_17853_),
    .B(_17857_),
    .Y(_17858_));
 sky130_fd_sc_hd__a21oi_2 _40234_ (.A1(_17702_),
    .A2(_17701_),
    .B1(_17682_),
    .Y(_17859_));
 sky130_fd_sc_hd__a21oi_1 _40235_ (.A1(_17726_),
    .A2(_17703_),
    .B1(_17859_),
    .Y(_17860_));
 sky130_fd_sc_hd__nand2_2 _40236_ (.A(_17858_),
    .B(_17860_),
    .Y(_17861_));
 sky130_fd_sc_hd__a21o_1 _40237_ (.A1(_17726_),
    .A2(_17703_),
    .B1(_17859_),
    .X(_17862_));
 sky130_fd_sc_hd__nand3_4 _40238_ (.A(_17862_),
    .B(_17857_),
    .C(_17853_),
    .Y(_17863_));
 sky130_fd_sc_hd__o21a_2 _40239_ (.A1(_16802_),
    .A2(_17249_),
    .B1(_17434_),
    .X(_17864_));
 sky130_fd_sc_hd__o21a_1 _40240_ (.A1(_17709_),
    .A2(_17720_),
    .B1(_17719_),
    .X(_17865_));
 sky130_fd_sc_hd__nor2_1 _40241_ (.A(_17864_),
    .B(_17865_),
    .Y(_17866_));
 sky130_fd_sc_hd__nand2_1 _40242_ (.A(_17865_),
    .B(_17864_),
    .Y(_17867_));
 sky130_fd_sc_hd__or2b_2 _40243_ (.A(_17866_),
    .B_N(_17867_),
    .X(_17868_));
 sky130_fd_sc_hd__a21oi_2 _40244_ (.A1(_17861_),
    .A2(_17863_),
    .B1(_17868_),
    .Y(_17869_));
 sky130_vsdinv _40245_ (.A(_17867_),
    .Y(_17870_));
 sky130_fd_sc_hd__o211a_1 _40246_ (.A1(_17870_),
    .A2(_17866_),
    .B1(_17863_),
    .C1(_17861_),
    .X(_17871_));
 sky130_fd_sc_hd__nand2_1 _40247_ (.A(_17679_),
    .B(_17675_),
    .Y(_17872_));
 sky130_fd_sc_hd__o22ai_4 _40248_ (.A1(_17732_),
    .A2(_17735_),
    .B1(_17872_),
    .B2(_17729_),
    .Y(_17873_));
 sky130_fd_sc_hd__o21bai_4 _40249_ (.A1(_17869_),
    .A2(_17871_),
    .B1_N(_17873_),
    .Y(_17874_));
 sky130_fd_sc_hd__a21o_1 _40250_ (.A1(_17861_),
    .A2(_17863_),
    .B1(_17868_),
    .X(_17875_));
 sky130_fd_sc_hd__nand3_4 _40251_ (.A(_17861_),
    .B(_17868_),
    .C(_17863_),
    .Y(_17876_));
 sky130_fd_sc_hd__nand3_4 _40252_ (.A(_17875_),
    .B(_17873_),
    .C(_17876_),
    .Y(_17877_));
 sky130_fd_sc_hd__a21o_1 _40253_ (.A1(_17675_),
    .A2(_17673_),
    .B1(_17167_),
    .X(_17878_));
 sky130_fd_sc_hd__nand3_2 _40254_ (.A(_17675_),
    .B(_17167_),
    .C(_17673_),
    .Y(_17879_));
 sky130_fd_sc_hd__a21o_1 _40255_ (.A1(_17878_),
    .A2(_17879_),
    .B1(_17613_),
    .X(_17880_));
 sky130_fd_sc_hd__nand3_1 _40256_ (.A(_17878_),
    .B(_17613_),
    .C(_17879_),
    .Y(_17881_));
 sky130_fd_sc_hd__nand2_2 _40257_ (.A(_17880_),
    .B(_17881_),
    .Y(_17882_));
 sky130_fd_sc_hd__a21o_1 _40258_ (.A1(_17874_),
    .A2(_17877_),
    .B1(_17882_),
    .X(_17883_));
 sky130_fd_sc_hd__o21ai_2 _40259_ (.A1(_17744_),
    .A2(_17741_),
    .B1(_17746_),
    .Y(_17884_));
 sky130_fd_sc_hd__nand3_4 _40260_ (.A(_17874_),
    .B(_17877_),
    .C(_17882_),
    .Y(_17885_));
 sky130_fd_sc_hd__nand3_4 _40261_ (.A(_17883_),
    .B(_17884_),
    .C(_17885_),
    .Y(_17886_));
 sky130_fd_sc_hd__a21oi_2 _40262_ (.A1(_17874_),
    .A2(_17877_),
    .B1(_17882_),
    .Y(_17887_));
 sky130_fd_sc_hd__nand2_1 _40263_ (.A(_17875_),
    .B(_17873_),
    .Y(_17888_));
 sky130_fd_sc_hd__o211a_1 _40264_ (.A1(_17871_),
    .A2(_17888_),
    .B1(_17882_),
    .C1(_17874_),
    .X(_17889_));
 sky130_fd_sc_hd__o21bai_4 _40265_ (.A1(_17887_),
    .A2(_17889_),
    .B1_N(_17884_),
    .Y(_17890_));
 sky130_fd_sc_hd__clkbuf_4 _40266_ (.A(_17476_),
    .X(_17891_));
 sky130_vsdinv _40267_ (.A(_17666_),
    .Y(_17892_));
 sky130_fd_sc_hd__a21o_1 _40268_ (.A1(_17665_),
    .A2(_17461_),
    .B1(_17892_),
    .X(_17893_));
 sky130_fd_sc_hd__nand2_1 _40269_ (.A(_17893_),
    .B(_17012_),
    .Y(_17894_));
 sky130_fd_sc_hd__clkbuf_4 _40270_ (.A(_17461_),
    .X(_17895_));
 sky130_fd_sc_hd__a211o_1 _40271_ (.A1(_17665_),
    .A2(_17895_),
    .B1(_17012_),
    .C1(_17892_),
    .X(_17896_));
 sky130_fd_sc_hd__nand2_1 _40272_ (.A(_17894_),
    .B(_17896_),
    .Y(_17897_));
 sky130_fd_sc_hd__nor2_1 _40273_ (.A(_17891_),
    .B(_17897_),
    .Y(_17898_));
 sky130_fd_sc_hd__and2_1 _40274_ (.A(_17897_),
    .B(_17476_),
    .X(_17899_));
 sky130_fd_sc_hd__o2bb2ai_2 _40275_ (.A1_N(_17886_),
    .A2_N(_17890_),
    .B1(_17898_),
    .B2(_17899_),
    .Y(_17900_));
 sky130_fd_sc_hd__nand2_1 _40276_ (.A(_17897_),
    .B(_17635_),
    .Y(_17901_));
 sky130_fd_sc_hd__nand3_1 _40277_ (.A(_17894_),
    .B(_17896_),
    .C(_17891_),
    .Y(_17902_));
 sky130_fd_sc_hd__nand2_2 _40278_ (.A(_17901_),
    .B(_17902_),
    .Y(_17903_));
 sky130_fd_sc_hd__nand3_4 _40279_ (.A(_17890_),
    .B(_17886_),
    .C(_17903_),
    .Y(_17904_));
 sky130_fd_sc_hd__o21ai_4 _40280_ (.A1(_17759_),
    .A2(_17750_),
    .B1(_17763_),
    .Y(_17905_));
 sky130_fd_sc_hd__a21oi_2 _40281_ (.A1(_17900_),
    .A2(_17904_),
    .B1(_17905_),
    .Y(_17906_));
 sky130_vsdinv _40282_ (.A(_17886_),
    .Y(_17907_));
 sky130_fd_sc_hd__nand2_1 _40283_ (.A(_17890_),
    .B(_17903_),
    .Y(_17908_));
 sky130_fd_sc_hd__o211a_2 _40284_ (.A1(_17907_),
    .A2(_17908_),
    .B1(_17905_),
    .C1(_17900_),
    .X(_17909_));
 sky130_fd_sc_hd__o22ai_4 _40285_ (.A1(_17808_),
    .A2(_17809_),
    .B1(_17906_),
    .B2(_17909_),
    .Y(_17910_));
 sky130_fd_sc_hd__a21o_1 _40286_ (.A1(_17900_),
    .A2(_17904_),
    .B1(_17905_),
    .X(_17911_));
 sky130_fd_sc_hd__nand3_2 _40287_ (.A(_17900_),
    .B(_17905_),
    .C(_17904_),
    .Y(_17912_));
 sky130_fd_sc_hd__nor2_2 _40288_ (.A(_17808_),
    .B(_17809_),
    .Y(_17913_));
 sky130_fd_sc_hd__nand3_4 _40289_ (.A(_17911_),
    .B(_17912_),
    .C(_17913_),
    .Y(_17914_));
 sky130_fd_sc_hd__o21ai_2 _40290_ (.A1(_17773_),
    .A2(_17767_),
    .B1(_17778_),
    .Y(_17915_));
 sky130_fd_sc_hd__a21oi_2 _40291_ (.A1(_17910_),
    .A2(_17914_),
    .B1(_17915_),
    .Y(_17916_));
 sky130_fd_sc_hd__a22oi_1 _40292_ (.A1(_17770_),
    .A2(_17771_),
    .B1(_17775_),
    .B2(_17776_),
    .Y(_17917_));
 sky130_fd_sc_hd__o211a_1 _40293_ (.A1(_17768_),
    .A2(_17917_),
    .B1(_17914_),
    .C1(_17910_),
    .X(_17918_));
 sky130_fd_sc_hd__o22ai_4 _40294_ (.A1(_17789_),
    .A2(_17769_),
    .B1(_17916_),
    .B2(_17918_),
    .Y(_17919_));
 sky130_fd_sc_hd__a21o_1 _40295_ (.A1(_17910_),
    .A2(_17914_),
    .B1(_17915_),
    .X(_17920_));
 sky130_fd_sc_hd__nor2_2 _40296_ (.A(_16515_),
    .B(_17769_),
    .Y(_17921_));
 sky130_fd_sc_hd__nand3_2 _40297_ (.A(_17915_),
    .B(_17910_),
    .C(_17914_),
    .Y(_17922_));
 sky130_fd_sc_hd__nand3_4 _40298_ (.A(_17920_),
    .B(_17921_),
    .C(_17922_),
    .Y(_17923_));
 sky130_fd_sc_hd__nand2_1 _40299_ (.A(_17786_),
    .B(_17662_),
    .Y(_17924_));
 sky130_fd_sc_hd__nand2_1 _40300_ (.A(_17924_),
    .B(_17782_),
    .Y(_17925_));
 sky130_fd_sc_hd__a21oi_4 _40301_ (.A1(_17919_),
    .A2(_17923_),
    .B1(_17925_),
    .Y(_17926_));
 sky130_fd_sc_hd__and3_1 _40302_ (.A(_17774_),
    .B(_17779_),
    .C(_17781_),
    .X(_17927_));
 sky130_fd_sc_hd__a31oi_1 _40303_ (.A1(_17783_),
    .A2(_17784_),
    .A3(_17785_),
    .B1(_17663_),
    .Y(_17928_));
 sky130_fd_sc_hd__o211a_2 _40304_ (.A1(_17927_),
    .A2(_17928_),
    .B1(_17923_),
    .C1(_17919_),
    .X(_17929_));
 sky130_fd_sc_hd__nor2_8 _40305_ (.A(_17926_),
    .B(_17929_),
    .Y(_17930_));
 sky130_fd_sc_hd__nor2_1 _40306_ (.A(_17788_),
    .B(_17793_),
    .Y(_17931_));
 sky130_fd_sc_hd__o21ai_2 _40307_ (.A1(_17931_),
    .A2(_17805_),
    .B1(_17796_),
    .Y(_17932_));
 sky130_fd_sc_hd__xnor2_2 _40308_ (.A(_17930_),
    .B(_17932_),
    .Y(_02678_));
 sky130_fd_sc_hd__a21o_1 _40309_ (.A1(_17920_),
    .A2(_17921_),
    .B1(_17918_),
    .X(_17933_));
 sky130_fd_sc_hd__and2_1 _40310_ (.A(_17857_),
    .B(_17842_),
    .X(_17934_));
 sky130_fd_sc_hd__nor2_1 _40311_ (.A(net465),
    .B(_15834_),
    .Y(_17935_));
 sky130_fd_sc_hd__a21oi_1 _40312_ (.A1(_19585_),
    .A2(_19828_),
    .B1(_17935_),
    .Y(_17936_));
 sky130_fd_sc_hd__and3_1 _40313_ (.A(_17935_),
    .B(_19585_),
    .C(_19828_),
    .X(_17937_));
 sky130_fd_sc_hd__nor2_1 _40314_ (.A(_17936_),
    .B(_17937_),
    .Y(_17938_));
 sky130_fd_sc_hd__or2_1 _40315_ (.A(_17829_),
    .B(_17938_),
    .X(_17939_));
 sky130_fd_sc_hd__nand2_1 _40316_ (.A(_17938_),
    .B(_17829_),
    .Y(_17940_));
 sky130_fd_sc_hd__nand2_1 _40317_ (.A(_17939_),
    .B(_17940_),
    .Y(_17941_));
 sky130_fd_sc_hd__nand2_1 _40318_ (.A(_19581_),
    .B(_19832_),
    .Y(_17942_));
 sky130_fd_sc_hd__or4_4 _40319_ (.A(_19841_),
    .B(_18476_),
    .C(_16353_),
    .D(_15780_),
    .X(_17943_));
 sky130_fd_sc_hd__a22o_1 _40320_ (.A1(_19578_),
    .A2(_19836_),
    .B1(_12902_),
    .B2(_11294_),
    .X(_17944_));
 sky130_fd_sc_hd__nand2_1 _40321_ (.A(_17943_),
    .B(_17944_),
    .Y(_17945_));
 sky130_fd_sc_hd__or2_2 _40322_ (.A(_17942_),
    .B(_17945_),
    .X(_17946_));
 sky130_fd_sc_hd__nand2_1 _40323_ (.A(_17945_),
    .B(_17942_),
    .Y(_17947_));
 sky130_fd_sc_hd__nand2_1 _40324_ (.A(_17946_),
    .B(_17947_),
    .Y(_17948_));
 sky130_fd_sc_hd__a21o_1 _40325_ (.A1(_17814_),
    .A2(_17818_),
    .B1(_17948_),
    .X(_17949_));
 sky130_fd_sc_hd__nand3_1 _40326_ (.A(_17948_),
    .B(_17814_),
    .C(_17818_),
    .Y(_17950_));
 sky130_fd_sc_hd__nand2_2 _40327_ (.A(_17949_),
    .B(_17950_),
    .Y(_17951_));
 sky130_fd_sc_hd__or2_1 _40328_ (.A(_17941_),
    .B(_17951_),
    .X(_17952_));
 sky130_fd_sc_hd__nand2_1 _40329_ (.A(_17840_),
    .B(_17820_),
    .Y(_17953_));
 sky130_fd_sc_hd__nand2_1 _40330_ (.A(_17951_),
    .B(_17941_),
    .Y(_17954_));
 sky130_fd_sc_hd__and3_1 _40331_ (.A(_17952_),
    .B(_17953_),
    .C(_17954_),
    .X(_17955_));
 sky130_vsdinv _40332_ (.A(_17941_),
    .Y(_17956_));
 sky130_fd_sc_hd__or2_1 _40333_ (.A(_17956_),
    .B(_17951_),
    .X(_17957_));
 sky130_vsdinv _40334_ (.A(_17953_),
    .Y(_17958_));
 sky130_fd_sc_hd__nand2_1 _40335_ (.A(_17951_),
    .B(_17956_),
    .Y(_17959_));
 sky130_fd_sc_hd__and3_1 _40336_ (.A(_17957_),
    .B(_17958_),
    .C(_17959_),
    .X(_17960_));
 sky130_fd_sc_hd__a21o_1 _40337_ (.A1(_17827_),
    .A2(_17829_),
    .B1(_17825_),
    .X(_17961_));
 sky130_fd_sc_hd__buf_1 _40338_ (.A(_17717_),
    .X(_17962_));
 sky130_fd_sc_hd__or2_1 _40339_ (.A(_17961_),
    .B(_17962_),
    .X(_17963_));
 sky130_fd_sc_hd__nand2_1 _40340_ (.A(_17962_),
    .B(_17961_),
    .Y(_17964_));
 sky130_fd_sc_hd__nand2_1 _40341_ (.A(_17963_),
    .B(_17964_),
    .Y(_17965_));
 sky130_fd_sc_hd__or2_2 _40342_ (.A(_17845_),
    .B(_17965_),
    .X(_17966_));
 sky130_fd_sc_hd__nand2_1 _40343_ (.A(_17965_),
    .B(_17846_),
    .Y(_17967_));
 sky130_fd_sc_hd__nand2_2 _40344_ (.A(_17966_),
    .B(_17967_),
    .Y(_17968_));
 sky130_fd_sc_hd__o21ai_2 _40345_ (.A1(_17955_),
    .A2(_17960_),
    .B1(_17968_),
    .Y(_17969_));
 sky130_fd_sc_hd__a21o_1 _40346_ (.A1(_17957_),
    .A2(_17959_),
    .B1(_17958_),
    .X(_17970_));
 sky130_fd_sc_hd__a21o_1 _40347_ (.A1(_17952_),
    .A2(_17954_),
    .B1(_17953_),
    .X(_17971_));
 sky130_vsdinv _40348_ (.A(_17968_),
    .Y(_17972_));
 sky130_fd_sc_hd__nand3_2 _40349_ (.A(_17970_),
    .B(_17971_),
    .C(_17972_),
    .Y(_17973_));
 sky130_fd_sc_hd__nand3b_4 _40350_ (.A_N(_17934_),
    .B(_17969_),
    .C(_17973_),
    .Y(_17974_));
 sky130_fd_sc_hd__o21ai_2 _40351_ (.A1(_17955_),
    .A2(_17960_),
    .B1(_17972_),
    .Y(_17975_));
 sky130_fd_sc_hd__nand3_2 _40352_ (.A(_17970_),
    .B(_17971_),
    .C(_17968_),
    .Y(_17976_));
 sky130_fd_sc_hd__nand3_4 _40353_ (.A(_17975_),
    .B(_17934_),
    .C(_17976_),
    .Y(_17977_));
 sky130_fd_sc_hd__o21ai_1 _40354_ (.A1(_17845_),
    .A2(_17850_),
    .B1(_17849_),
    .Y(_17978_));
 sky130_fd_sc_hd__or2_1 _40355_ (.A(_17586_),
    .B(_17978_),
    .X(_17979_));
 sky130_fd_sc_hd__nand2_1 _40356_ (.A(_17978_),
    .B(_17586_),
    .Y(_17980_));
 sky130_fd_sc_hd__nand2_2 _40357_ (.A(_17979_),
    .B(_17980_),
    .Y(_17981_));
 sky130_fd_sc_hd__xor2_4 _40358_ (.A(_17591_),
    .B(_17981_),
    .X(_17982_));
 sky130_fd_sc_hd__a21oi_4 _40359_ (.A1(_17974_),
    .A2(_17977_),
    .B1(_17982_),
    .Y(_17983_));
 sky130_fd_sc_hd__and3_1 _40360_ (.A(_17974_),
    .B(_17977_),
    .C(_17982_),
    .X(_17984_));
 sky130_fd_sc_hd__nand2_2 _40361_ (.A(_17876_),
    .B(_17863_),
    .Y(_17985_));
 sky130_fd_sc_hd__o21bai_4 _40362_ (.A1(_17983_),
    .A2(_17984_),
    .B1_N(_17985_),
    .Y(_17986_));
 sky130_fd_sc_hd__nand3_4 _40363_ (.A(_17974_),
    .B(_17977_),
    .C(_17982_),
    .Y(_17987_));
 sky130_fd_sc_hd__nand3b_4 _40364_ (.A_N(_17983_),
    .B(_17985_),
    .C(_17987_),
    .Y(_17988_));
 sky130_fd_sc_hd__o21ai_2 _40365_ (.A1(_17436_),
    .A2(_17865_),
    .B1(_17434_),
    .Y(_17989_));
 sky130_fd_sc_hd__nor2_2 _40366_ (.A(_17607_),
    .B(_17989_),
    .Y(_17990_));
 sky130_fd_sc_hd__and2_1 _40367_ (.A(_17989_),
    .B(_17607_),
    .X(_17991_));
 sky130_fd_sc_hd__nor2_4 _40368_ (.A(_17990_),
    .B(_17991_),
    .Y(_17992_));
 sky130_fd_sc_hd__xor2_4 _40369_ (.A(_17895_),
    .B(_17992_),
    .X(_17993_));
 sky130_fd_sc_hd__a21oi_1 _40370_ (.A1(_17986_),
    .A2(_17988_),
    .B1(_17993_),
    .Y(_17994_));
 sky130_fd_sc_hd__and3_1 _40371_ (.A(_17986_),
    .B(_17988_),
    .C(_17993_),
    .X(_17995_));
 sky130_fd_sc_hd__nand2_2 _40372_ (.A(_17885_),
    .B(_17877_),
    .Y(_17996_));
 sky130_fd_sc_hd__o21bai_2 _40373_ (.A1(_17994_),
    .A2(_17995_),
    .B1_N(_17996_),
    .Y(_17997_));
 sky130_fd_sc_hd__a21o_1 _40374_ (.A1(_17986_),
    .A2(_17988_),
    .B1(_17993_),
    .X(_17998_));
 sky130_fd_sc_hd__nand3_4 _40375_ (.A(_17986_),
    .B(_17988_),
    .C(_17993_),
    .Y(_17999_));
 sky130_fd_sc_hd__nand3_4 _40376_ (.A(_17998_),
    .B(_17996_),
    .C(_17999_),
    .Y(_18000_));
 sky130_fd_sc_hd__nand2_1 _40377_ (.A(_17997_),
    .B(_18000_),
    .Y(_18001_));
 sky130_fd_sc_hd__clkbuf_2 _40378_ (.A(_17012_),
    .X(_18002_));
 sky130_fd_sc_hd__a21bo_1 _40379_ (.A1(_17461_),
    .A2(_17879_),
    .B1_N(_17878_),
    .X(_18003_));
 sky130_fd_sc_hd__or2_1 _40380_ (.A(_18002_),
    .B(_18003_),
    .X(_18004_));
 sky130_fd_sc_hd__nand2_1 _40381_ (.A(_18003_),
    .B(_18002_),
    .Y(_18005_));
 sky130_fd_sc_hd__nand2_2 _40382_ (.A(_18004_),
    .B(_18005_),
    .Y(_18006_));
 sky130_fd_sc_hd__nor2_2 _40383_ (.A(_17806_),
    .B(_18006_),
    .Y(_18007_));
 sky130_fd_sc_hd__and2_1 _40384_ (.A(_18006_),
    .B(_17635_),
    .X(_18008_));
 sky130_fd_sc_hd__nor2_4 _40385_ (.A(_18007_),
    .B(_18008_),
    .Y(_18009_));
 sky130_fd_sc_hd__nand2_1 _40386_ (.A(_18001_),
    .B(_18009_),
    .Y(_18010_));
 sky130_fd_sc_hd__nand2_2 _40387_ (.A(_17908_),
    .B(_17886_),
    .Y(_18011_));
 sky130_vsdinv _40388_ (.A(_18009_),
    .Y(_18012_));
 sky130_fd_sc_hd__nand3_2 _40389_ (.A(_18012_),
    .B(_17997_),
    .C(_18000_),
    .Y(_18013_));
 sky130_fd_sc_hd__nand3_4 _40390_ (.A(_18010_),
    .B(_18011_),
    .C(_18013_),
    .Y(_18014_));
 sky130_fd_sc_hd__nand2_1 _40391_ (.A(_18001_),
    .B(_18012_),
    .Y(_18015_));
 sky130_vsdinv _40392_ (.A(_18011_),
    .Y(_18016_));
 sky130_fd_sc_hd__nand3_2 _40393_ (.A(_17997_),
    .B(_18000_),
    .C(_18009_),
    .Y(_18017_));
 sky130_fd_sc_hd__nand3_4 _40394_ (.A(_18015_),
    .B(_18016_),
    .C(_18017_),
    .Y(_18018_));
 sky130_fd_sc_hd__nand2_1 _40395_ (.A(_17896_),
    .B(_17806_),
    .Y(_18019_));
 sky130_fd_sc_hd__nand2_2 _40396_ (.A(_18019_),
    .B(_17894_),
    .Y(_18020_));
 sky130_fd_sc_hd__nor2_4 _40397_ (.A(_16515_),
    .B(_18020_),
    .Y(_18021_));
 sky130_vsdinv _40398_ (.A(_18020_),
    .Y(_18022_));
 sky130_fd_sc_hd__nor2_4 _40399_ (.A(_17353_),
    .B(_18022_),
    .Y(_18023_));
 sky130_fd_sc_hd__nor2_2 _40400_ (.A(_18021_),
    .B(_18023_),
    .Y(_18024_));
 sky130_fd_sc_hd__nand3_4 _40401_ (.A(_18014_),
    .B(_18018_),
    .C(_18024_),
    .Y(_18025_));
 sky130_fd_sc_hd__o2bb2ai_2 _40402_ (.A1_N(_18018_),
    .A2_N(_18014_),
    .B1(_18021_),
    .B2(_18023_),
    .Y(_18026_));
 sky130_vsdinv _40403_ (.A(_17914_),
    .Y(_18027_));
 sky130_fd_sc_hd__o2bb2ai_2 _40404_ (.A1_N(_18025_),
    .A2_N(_18026_),
    .B1(_17909_),
    .B2(_18027_),
    .Y(_18028_));
 sky130_fd_sc_hd__nor2_2 _40405_ (.A(_17909_),
    .B(_18027_),
    .Y(_18029_));
 sky130_fd_sc_hd__nand3_4 _40406_ (.A(_18026_),
    .B(_18029_),
    .C(_18025_),
    .Y(_18030_));
 sky130_fd_sc_hd__nand2_1 _40407_ (.A(_18028_),
    .B(_18030_),
    .Y(_18031_));
 sky130_fd_sc_hd__nand2_1 _40408_ (.A(_18031_),
    .B(_17808_),
    .Y(_18032_));
 sky130_vsdinv _40409_ (.A(_17808_),
    .Y(_18033_));
 sky130_fd_sc_hd__nand3_2 _40410_ (.A(_18028_),
    .B(_18033_),
    .C(_18030_),
    .Y(_18034_));
 sky130_fd_sc_hd__nand3b_4 _40411_ (.A_N(_17933_),
    .B(_18032_),
    .C(_18034_),
    .Y(_18035_));
 sky130_fd_sc_hd__nand2_1 _40412_ (.A(_18031_),
    .B(_18033_),
    .Y(_18036_));
 sky130_fd_sc_hd__nand3_2 _40413_ (.A(_18028_),
    .B(_17808_),
    .C(_18030_),
    .Y(_18037_));
 sky130_fd_sc_hd__nand3_4 _40414_ (.A(_18036_),
    .B(_17933_),
    .C(_18037_),
    .Y(_18038_));
 sky130_fd_sc_hd__nand2_2 _40415_ (.A(_18035_),
    .B(_18038_),
    .Y(_18039_));
 sky130_fd_sc_hd__nand3_1 _40416_ (.A(_17801_),
    .B(_17930_),
    .C(_17797_),
    .Y(_18040_));
 sky130_fd_sc_hd__o21bai_4 _40417_ (.A1(_17518_),
    .A2(_17522_),
    .B1_N(_18040_),
    .Y(_18041_));
 sky130_vsdinv _40418_ (.A(_17929_),
    .Y(_18042_));
 sky130_fd_sc_hd__o31ai_4 _40419_ (.A1(_17788_),
    .A2(_17793_),
    .A3(_17926_),
    .B1(_18042_),
    .Y(_18043_));
 sky130_fd_sc_hd__a31oi_4 _40420_ (.A1(_17804_),
    .A2(_17797_),
    .A3(_17930_),
    .B1(_18043_),
    .Y(_18044_));
 sky130_fd_sc_hd__nand2_4 _40421_ (.A(_18041_),
    .B(_18044_),
    .Y(_18045_));
 sky130_fd_sc_hd__xnor2_4 _40422_ (.A(_18039_),
    .B(_18045_),
    .Y(_02679_));
 sky130_fd_sc_hd__a21o_1 _40423_ (.A1(_17992_),
    .A2(_17895_),
    .B1(_17991_),
    .X(_18046_));
 sky130_fd_sc_hd__or2_1 _40424_ (.A(_18002_),
    .B(_18046_),
    .X(_18047_));
 sky130_fd_sc_hd__nand2_1 _40425_ (.A(_18046_),
    .B(_18002_),
    .Y(_18048_));
 sky130_fd_sc_hd__nand2_2 _40426_ (.A(_18047_),
    .B(_18048_),
    .Y(_18049_));
 sky130_fd_sc_hd__nor2_8 _40427_ (.A(_17891_),
    .B(_18049_),
    .Y(_18050_));
 sky130_fd_sc_hd__and2_2 _40428_ (.A(_18049_),
    .B(_17891_),
    .X(_18051_));
 sky130_fd_sc_hd__o21ai_2 _40429_ (.A1(_17968_),
    .A2(_17960_),
    .B1(_17970_),
    .Y(_18052_));
 sky130_fd_sc_hd__or4_4 _40430_ (.A(_19836_),
    .B(_18476_),
    .C(_16353_),
    .D(_17288_),
    .X(_18053_));
 sky130_fd_sc_hd__a22o_1 _40431_ (.A1(_19578_),
    .A2(_19832_),
    .B1(_15780_),
    .B2(_11294_),
    .X(_18054_));
 sky130_fd_sc_hd__nand2_1 _40432_ (.A(_18053_),
    .B(_18054_),
    .Y(_18055_));
 sky130_fd_sc_hd__or3_1 _40433_ (.A(_15814_),
    .B(_17245_),
    .C(_18055_),
    .X(_18056_));
 sky130_fd_sc_hd__o21ai_1 _40434_ (.A1(_15814_),
    .A2(_17245_),
    .B1(_18055_),
    .Y(_18057_));
 sky130_fd_sc_hd__nand2_2 _40435_ (.A(_18056_),
    .B(_18057_),
    .Y(_18058_));
 sky130_fd_sc_hd__a21o_2 _40436_ (.A1(_17943_),
    .A2(_17946_),
    .B1(_18058_),
    .X(_18059_));
 sky130_fd_sc_hd__nand3_4 _40437_ (.A(_18058_),
    .B(_17943_),
    .C(_17946_),
    .Y(_18060_));
 sky130_fd_sc_hd__o21ai_1 _40438_ (.A1(_19585_),
    .A2(_19589_),
    .B1(_14218_),
    .Y(_18061_));
 sky130_fd_sc_hd__and3_1 _40439_ (.A(_14218_),
    .B(_19585_),
    .C(_19589_),
    .X(_18062_));
 sky130_fd_sc_hd__nor2_2 _40440_ (.A(_18061_),
    .B(_18062_),
    .Y(_18063_));
 sky130_fd_sc_hd__nor2_4 _40441_ (.A(_17829_),
    .B(_18063_),
    .Y(_18064_));
 sky130_fd_sc_hd__and2_2 _40442_ (.A(_18063_),
    .B(_19594_),
    .X(_18065_));
 sky130_fd_sc_hd__nor2_8 _40443_ (.A(_18064_),
    .B(_18065_),
    .Y(_18066_));
 sky130_fd_sc_hd__a21o_1 _40444_ (.A1(_18059_),
    .A2(_18060_),
    .B1(_18066_),
    .X(_18067_));
 sky130_fd_sc_hd__nand3_4 _40445_ (.A(_18059_),
    .B(_18066_),
    .C(_18060_),
    .Y(_18068_));
 sky130_fd_sc_hd__o21a_1 _40446_ (.A1(_17941_),
    .A2(_17951_),
    .B1(_17949_),
    .X(_18069_));
 sky130_fd_sc_hd__a21bo_1 _40447_ (.A1(_18067_),
    .A2(_18068_),
    .B1_N(_18069_),
    .X(_18070_));
 sky130_fd_sc_hd__nand3b_4 _40448_ (.A_N(_18069_),
    .B(_18068_),
    .C(_18067_),
    .Y(_18071_));
 sky130_fd_sc_hd__nand2_1 _40449_ (.A(_18070_),
    .B(_18071_),
    .Y(_18072_));
 sky130_fd_sc_hd__a21o_1 _40450_ (.A1(_17938_),
    .A2(_17829_),
    .B1(_17937_),
    .X(_18073_));
 sky130_fd_sc_hd__or2_1 _40451_ (.A(_18073_),
    .B(_17962_),
    .X(_18074_));
 sky130_fd_sc_hd__nand2_1 _40452_ (.A(_17962_),
    .B(_18073_),
    .Y(_18075_));
 sky130_fd_sc_hd__nand2_1 _40453_ (.A(_18074_),
    .B(_18075_),
    .Y(_18076_));
 sky130_fd_sc_hd__or2_1 _40454_ (.A(_17845_),
    .B(_18076_),
    .X(_18077_));
 sky130_fd_sc_hd__nand2_1 _40455_ (.A(_18076_),
    .B(_17846_),
    .Y(_18078_));
 sky130_fd_sc_hd__nand2_1 _40456_ (.A(_18077_),
    .B(_18078_),
    .Y(_18079_));
 sky130_vsdinv _40457_ (.A(_18079_),
    .Y(_18080_));
 sky130_fd_sc_hd__nand2_1 _40458_ (.A(_18072_),
    .B(_18080_),
    .Y(_18081_));
 sky130_fd_sc_hd__nand3_2 _40459_ (.A(_18070_),
    .B(_18079_),
    .C(_18071_),
    .Y(_18082_));
 sky130_fd_sc_hd__nand3b_4 _40460_ (.A_N(_18052_),
    .B(_18081_),
    .C(_18082_),
    .Y(_18083_));
 sky130_fd_sc_hd__nand2_1 _40461_ (.A(_18072_),
    .B(_18079_),
    .Y(_18084_));
 sky130_fd_sc_hd__nand3_4 _40462_ (.A(_18070_),
    .B(_18080_),
    .C(_18071_),
    .Y(_18085_));
 sky130_fd_sc_hd__nand3_4 _40463_ (.A(_18084_),
    .B(_18052_),
    .C(_18085_),
    .Y(_18086_));
 sky130_fd_sc_hd__nand2_1 _40464_ (.A(_17966_),
    .B(_17964_),
    .Y(_18087_));
 sky130_fd_sc_hd__nand2_1 _40465_ (.A(_18087_),
    .B(_17586_),
    .Y(_18088_));
 sky130_fd_sc_hd__nand3_2 _40466_ (.A(_17966_),
    .B(_17588_),
    .C(_17964_),
    .Y(_18089_));
 sky130_fd_sc_hd__a21oi_2 _40467_ (.A1(_18088_),
    .A2(_18089_),
    .B1(_17585_),
    .Y(_18090_));
 sky130_fd_sc_hd__and3_1 _40468_ (.A(_18088_),
    .B(_17585_),
    .C(_18089_),
    .X(_18091_));
 sky130_fd_sc_hd__nor2_4 _40469_ (.A(_18090_),
    .B(_18091_),
    .Y(_18092_));
 sky130_fd_sc_hd__a21oi_4 _40470_ (.A1(_18083_),
    .A2(_18086_),
    .B1(_18092_),
    .Y(_18093_));
 sky130_fd_sc_hd__and3_1 _40471_ (.A(_18083_),
    .B(_18086_),
    .C(_18092_),
    .X(_18094_));
 sky130_fd_sc_hd__nand2_2 _40472_ (.A(_17987_),
    .B(_17974_),
    .Y(_18095_));
 sky130_fd_sc_hd__o21bai_4 _40473_ (.A1(_18093_),
    .A2(_18094_),
    .B1_N(_18095_),
    .Y(_18096_));
 sky130_fd_sc_hd__nand3_4 _40474_ (.A(_18083_),
    .B(_18086_),
    .C(_18092_),
    .Y(_18097_));
 sky130_fd_sc_hd__nand3b_4 _40475_ (.A_N(_18093_),
    .B(_18095_),
    .C(_18097_),
    .Y(_18098_));
 sky130_fd_sc_hd__o21a_1 _40476_ (.A1(_17591_),
    .A2(_17981_),
    .B1(_17980_),
    .X(_18099_));
 sky130_fd_sc_hd__or2_1 _40477_ (.A(_17167_),
    .B(_18099_),
    .X(_18100_));
 sky130_fd_sc_hd__nand2_1 _40478_ (.A(_18099_),
    .B(_17167_),
    .Y(_18101_));
 sky130_fd_sc_hd__a21o_1 _40479_ (.A1(_18100_),
    .A2(_18101_),
    .B1(_17613_),
    .X(_18102_));
 sky130_fd_sc_hd__nand3_1 _40480_ (.A(_18100_),
    .B(_17613_),
    .C(_18101_),
    .Y(_18103_));
 sky130_fd_sc_hd__nand2_2 _40481_ (.A(_18102_),
    .B(_18103_),
    .Y(_18104_));
 sky130_fd_sc_hd__a21o_2 _40482_ (.A1(_18096_),
    .A2(_18098_),
    .B1(_18104_),
    .X(_18105_));
 sky130_fd_sc_hd__nand3_4 _40483_ (.A(_18096_),
    .B(_18098_),
    .C(_18104_),
    .Y(_18106_));
 sky130_fd_sc_hd__nand2_2 _40484_ (.A(_17999_),
    .B(_17988_),
    .Y(_18107_));
 sky130_fd_sc_hd__a21oi_4 _40485_ (.A1(_18105_),
    .A2(_18106_),
    .B1(_18107_),
    .Y(_18108_));
 sky130_fd_sc_hd__a21boi_2 _40486_ (.A1(_17986_),
    .A2(_17993_),
    .B1_N(_17988_),
    .Y(_18109_));
 sky130_fd_sc_hd__a21oi_2 _40487_ (.A1(_18096_),
    .A2(_18098_),
    .B1(_18104_),
    .Y(_18110_));
 sky130_fd_sc_hd__nor3b_4 _40488_ (.A(_18109_),
    .B(_18110_),
    .C_N(_18106_),
    .Y(_18111_));
 sky130_fd_sc_hd__o22ai_4 _40489_ (.A1(_18050_),
    .A2(_18051_),
    .B1(_18108_),
    .B2(_18111_),
    .Y(_18112_));
 sky130_fd_sc_hd__a21oi_2 _40490_ (.A1(_17998_),
    .A2(_17999_),
    .B1(_17996_),
    .Y(_18113_));
 sky130_fd_sc_hd__o21ai_2 _40491_ (.A1(_18009_),
    .A2(_18113_),
    .B1(_18000_),
    .Y(_18114_));
 sky130_fd_sc_hd__a21o_1 _40492_ (.A1(_18105_),
    .A2(_18106_),
    .B1(_18107_),
    .X(_18115_));
 sky130_fd_sc_hd__nand3_4 _40493_ (.A(_18105_),
    .B(_18107_),
    .C(_18106_),
    .Y(_18116_));
 sky130_fd_sc_hd__nor2_8 _40494_ (.A(_18050_),
    .B(_18051_),
    .Y(_18117_));
 sky130_fd_sc_hd__nand3_4 _40495_ (.A(_18115_),
    .B(_18116_),
    .C(_18117_),
    .Y(_18118_));
 sky130_fd_sc_hd__nand3_4 _40496_ (.A(_18112_),
    .B(_18114_),
    .C(_18118_),
    .Y(_18119_));
 sky130_fd_sc_hd__o21ai_2 _40497_ (.A1(_18108_),
    .A2(_18111_),
    .B1(_18117_),
    .Y(_18120_));
 sky130_fd_sc_hd__o21a_1 _40498_ (.A1(_18009_),
    .A2(_18113_),
    .B1(_18000_),
    .X(_18121_));
 sky130_fd_sc_hd__nand3b_4 _40499_ (.A_N(_18117_),
    .B(_18115_),
    .C(_18116_),
    .Y(_18122_));
 sky130_fd_sc_hd__nand3_4 _40500_ (.A(_18120_),
    .B(_18121_),
    .C(_18122_),
    .Y(_18123_));
 sky130_fd_sc_hd__o21ai_2 _40501_ (.A1(_17891_),
    .A2(_18006_),
    .B1(_18005_),
    .Y(_18124_));
 sky130_fd_sc_hd__and2_2 _40502_ (.A(_18124_),
    .B(_17353_),
    .X(_18125_));
 sky130_fd_sc_hd__nor2_4 _40503_ (.A(_17353_),
    .B(_18124_),
    .Y(_18126_));
 sky130_fd_sc_hd__o2bb2ai_4 _40504_ (.A1_N(_18119_),
    .A2_N(_18123_),
    .B1(_18125_),
    .B2(_18126_),
    .Y(_18127_));
 sky130_fd_sc_hd__nor2_2 _40505_ (.A(_18126_),
    .B(_18125_),
    .Y(_18128_));
 sky130_fd_sc_hd__nand3_4 _40506_ (.A(_18123_),
    .B(_18119_),
    .C(_18128_),
    .Y(_18129_));
 sky130_fd_sc_hd__o21ai_2 _40507_ (.A1(_18021_),
    .A2(_18023_),
    .B1(_18018_),
    .Y(_18130_));
 sky130_fd_sc_hd__nand2_4 _40508_ (.A(_18130_),
    .B(_18014_),
    .Y(_18131_));
 sky130_fd_sc_hd__a21oi_4 _40509_ (.A1(_18127_),
    .A2(_18129_),
    .B1(_18131_),
    .Y(_18132_));
 sky130_fd_sc_hd__and3_1 _40510_ (.A(_18112_),
    .B(_18114_),
    .C(_18118_),
    .X(_18133_));
 sky130_fd_sc_hd__nand2_1 _40511_ (.A(_18123_),
    .B(_18128_),
    .Y(_18134_));
 sky130_fd_sc_hd__o211a_2 _40512_ (.A1(_18133_),
    .A2(_18134_),
    .B1(_18131_),
    .C1(_18127_),
    .X(_18135_));
 sky130_fd_sc_hd__nor2_1 _40513_ (.A(_17789_),
    .B(_18022_),
    .Y(_18136_));
 sky130_fd_sc_hd__o21ai_2 _40514_ (.A1(_18132_),
    .A2(_18135_),
    .B1(_18136_),
    .Y(_18137_));
 sky130_fd_sc_hd__nand3_4 _40515_ (.A(_18127_),
    .B(_18131_),
    .C(_18129_),
    .Y(_18138_));
 sky130_vsdinv _40516_ (.A(_18136_),
    .Y(_18139_));
 sky130_fd_sc_hd__nand3b_4 _40517_ (.A_N(_18132_),
    .B(_18138_),
    .C(_18139_),
    .Y(_18140_));
 sky130_fd_sc_hd__nand2_1 _40518_ (.A(_18030_),
    .B(_17808_),
    .Y(_18141_));
 sky130_fd_sc_hd__nand2_1 _40519_ (.A(_18141_),
    .B(_18028_),
    .Y(_18142_));
 sky130_fd_sc_hd__a21bo_1 _40520_ (.A1(_18137_),
    .A2(_18140_),
    .B1_N(_18142_),
    .X(_18143_));
 sky130_fd_sc_hd__nand3b_4 _40521_ (.A_N(_18142_),
    .B(_18137_),
    .C(_18140_),
    .Y(_18144_));
 sky130_fd_sc_hd__nand2_2 _40522_ (.A(_18143_),
    .B(_18144_),
    .Y(_18145_));
 sky130_vsdinv _40523_ (.A(_18038_),
    .Y(_18146_));
 sky130_fd_sc_hd__a21oi_4 _40524_ (.A1(_18045_),
    .A2(_18035_),
    .B1(_18146_),
    .Y(_18147_));
 sky130_fd_sc_hd__xor2_4 _40525_ (.A(_18145_),
    .B(_18147_),
    .X(_02680_));
 sky130_fd_sc_hd__nor2_4 _40526_ (.A(_18117_),
    .B(_18111_),
    .Y(_18148_));
 sky130_fd_sc_hd__and2_1 _40527_ (.A(_18097_),
    .B(_18086_),
    .X(_18149_));
 sky130_fd_sc_hd__nand2_2 _40528_ (.A(_18085_),
    .B(_18071_),
    .Y(_18150_));
 sky130_fd_sc_hd__nand2_2 _40529_ (.A(_18068_),
    .B(_18059_),
    .Y(_18151_));
 sky130_vsdinv _40530_ (.A(_18066_),
    .Y(_18152_));
 sky130_fd_sc_hd__nand2_4 _40531_ (.A(_14218_),
    .B(_19581_),
    .Y(_18153_));
 sky130_fd_sc_hd__and4_2 _40532_ (.A(_17288_),
    .B(_11294_),
    .C(_19578_),
    .D(_19828_),
    .X(_18154_));
 sky130_fd_sc_hd__o22a_1 _40533_ (.A1(_19832_),
    .A2(_18476_),
    .B1(_16353_),
    .B2(_17245_),
    .X(_18155_));
 sky130_fd_sc_hd__nor3_4 _40534_ (.A(_18153_),
    .B(_18154_),
    .C(_18155_),
    .Y(_18156_));
 sky130_fd_sc_hd__o21a_1 _40535_ (.A1(_18154_),
    .A2(_18155_),
    .B1(_18153_),
    .X(_18157_));
 sky130_fd_sc_hd__nor2_1 _40536_ (.A(_18156_),
    .B(_18157_),
    .Y(_18158_));
 sky130_fd_sc_hd__nand2_1 _40537_ (.A(_18056_),
    .B(_18053_),
    .Y(_18159_));
 sky130_fd_sc_hd__or2_1 _40538_ (.A(_18158_),
    .B(_18159_),
    .X(_18160_));
 sky130_fd_sc_hd__nand2_2 _40539_ (.A(_18159_),
    .B(_18158_),
    .Y(_18161_));
 sky130_fd_sc_hd__nand2_4 _40540_ (.A(_18160_),
    .B(_18161_),
    .Y(_18162_));
 sky130_fd_sc_hd__xor2_4 _40541_ (.A(_18152_),
    .B(_18162_),
    .X(_18163_));
 sky130_fd_sc_hd__or2_2 _40542_ (.A(_18151_),
    .B(_18163_),
    .X(_18164_));
 sky130_fd_sc_hd__nand2_4 _40543_ (.A(_18163_),
    .B(_18151_),
    .Y(_18165_));
 sky130_fd_sc_hd__nand2_1 _40544_ (.A(_18164_),
    .B(_18165_),
    .Y(_18166_));
 sky130_fd_sc_hd__or2_1 _40545_ (.A(_18062_),
    .B(_18065_),
    .X(_18167_));
 sky130_fd_sc_hd__or2_1 _40546_ (.A(_18167_),
    .B(_17962_),
    .X(_18168_));
 sky130_fd_sc_hd__nand2_1 _40547_ (.A(_17962_),
    .B(_18167_),
    .Y(_18169_));
 sky130_fd_sc_hd__nand2_1 _40548_ (.A(_18168_),
    .B(_18169_),
    .Y(_18170_));
 sky130_fd_sc_hd__or2_2 _40549_ (.A(_17846_),
    .B(_18170_),
    .X(_18171_));
 sky130_fd_sc_hd__nand2_1 _40550_ (.A(_18170_),
    .B(_17846_),
    .Y(_18172_));
 sky130_fd_sc_hd__nand2_4 _40551_ (.A(_18171_),
    .B(_18172_),
    .Y(_18173_));
 sky130_vsdinv _40552_ (.A(_18173_),
    .Y(_18174_));
 sky130_fd_sc_hd__nand2_1 _40553_ (.A(_18166_),
    .B(_18174_),
    .Y(_18175_));
 sky130_fd_sc_hd__nand3_2 _40554_ (.A(_18164_),
    .B(_18173_),
    .C(_18165_),
    .Y(_18176_));
 sky130_fd_sc_hd__nand3b_4 _40555_ (.A_N(_18150_),
    .B(_18175_),
    .C(_18176_),
    .Y(_18177_));
 sky130_fd_sc_hd__nand2_1 _40556_ (.A(_18166_),
    .B(_18173_),
    .Y(_18178_));
 sky130_fd_sc_hd__nand3_4 _40557_ (.A(_18164_),
    .B(_18174_),
    .C(_18165_),
    .Y(_18179_));
 sky130_fd_sc_hd__nand3_4 _40558_ (.A(_18178_),
    .B(_18150_),
    .C(_18179_),
    .Y(_18180_));
 sky130_fd_sc_hd__nand2_1 _40559_ (.A(_18177_),
    .B(_18180_),
    .Y(_18181_));
 sky130_fd_sc_hd__nand2_2 _40560_ (.A(_18077_),
    .B(_18075_),
    .Y(_18182_));
 sky130_fd_sc_hd__xnor2_2 _40561_ (.A(_17864_),
    .B(_18182_),
    .Y(_18183_));
 sky130_fd_sc_hd__nand2_1 _40562_ (.A(_18181_),
    .B(_18183_),
    .Y(_18184_));
 sky130_vsdinv _40563_ (.A(_18183_),
    .Y(_18185_));
 sky130_fd_sc_hd__nand3_4 _40564_ (.A(_18177_),
    .B(_18180_),
    .C(_18185_),
    .Y(_18186_));
 sky130_fd_sc_hd__nand3b_4 _40565_ (.A_N(_18149_),
    .B(_18184_),
    .C(_18186_),
    .Y(_18187_));
 sky130_fd_sc_hd__nand2_1 _40566_ (.A(_18181_),
    .B(_18185_),
    .Y(_18188_));
 sky130_fd_sc_hd__nand3_2 _40567_ (.A(_18177_),
    .B(_18180_),
    .C(_18183_),
    .Y(_18189_));
 sky130_fd_sc_hd__nand3_4 _40568_ (.A(_18188_),
    .B(_18189_),
    .C(_18149_),
    .Y(_18190_));
 sky130_vsdinv _40569_ (.A(_18088_),
    .Y(_18191_));
 sky130_fd_sc_hd__nor2_2 _40570_ (.A(_18191_),
    .B(_18091_),
    .Y(_18192_));
 sky130_fd_sc_hd__xor2_1 _40571_ (.A(_17607_),
    .B(_18192_),
    .X(_18193_));
 sky130_fd_sc_hd__nor2_1 _40572_ (.A(_17895_),
    .B(_18193_),
    .Y(_18194_));
 sky130_fd_sc_hd__nand2_1 _40573_ (.A(_18193_),
    .B(_17895_),
    .Y(_18195_));
 sky130_fd_sc_hd__or2b_2 _40574_ (.A(_18194_),
    .B_N(_18195_),
    .X(_18196_));
 sky130_fd_sc_hd__a21oi_2 _40575_ (.A1(_18187_),
    .A2(_18190_),
    .B1(_18196_),
    .Y(_18197_));
 sky130_vsdinv _40576_ (.A(_18195_),
    .Y(_18198_));
 sky130_fd_sc_hd__o211a_1 _40577_ (.A1(_18194_),
    .A2(_18198_),
    .B1(_18190_),
    .C1(_18187_),
    .X(_18199_));
 sky130_fd_sc_hd__nand2_2 _40578_ (.A(_18106_),
    .B(_18098_),
    .Y(_18200_));
 sky130_fd_sc_hd__o21bai_4 _40579_ (.A1(_18197_),
    .A2(_18199_),
    .B1_N(_18200_),
    .Y(_18201_));
 sky130_fd_sc_hd__a21o_1 _40580_ (.A1(_18187_),
    .A2(_18190_),
    .B1(_18196_),
    .X(_18202_));
 sky130_fd_sc_hd__nand3_2 _40581_ (.A(_18187_),
    .B(_18196_),
    .C(_18190_),
    .Y(_18203_));
 sky130_fd_sc_hd__nand3_4 _40582_ (.A(_18202_),
    .B(_18200_),
    .C(_18203_),
    .Y(_18204_));
 sky130_fd_sc_hd__nand2_1 _40583_ (.A(_18101_),
    .B(_17895_),
    .Y(_18205_));
 sky130_fd_sc_hd__nand2_1 _40584_ (.A(_18100_),
    .B(_18205_),
    .Y(_18206_));
 sky130_fd_sc_hd__or2_1 _40585_ (.A(_18002_),
    .B(_18206_),
    .X(_18207_));
 sky130_fd_sc_hd__nand2_1 _40586_ (.A(_18206_),
    .B(_18002_),
    .Y(_18208_));
 sky130_fd_sc_hd__nand2_1 _40587_ (.A(_18207_),
    .B(_18208_),
    .Y(_18209_));
 sky130_fd_sc_hd__nor2_1 _40588_ (.A(_17806_),
    .B(_18209_),
    .Y(_18210_));
 sky130_fd_sc_hd__and2_1 _40589_ (.A(_18209_),
    .B(_17806_),
    .X(_18211_));
 sky130_fd_sc_hd__or2_2 _40590_ (.A(_18210_),
    .B(_18211_),
    .X(_18212_));
 sky130_fd_sc_hd__a21oi_2 _40591_ (.A1(_18201_),
    .A2(_18204_),
    .B1(_18212_),
    .Y(_18213_));
 sky130_fd_sc_hd__o211a_1 _40592_ (.A1(_18211_),
    .A2(_18210_),
    .B1(_18204_),
    .C1(_18201_),
    .X(_18214_));
 sky130_fd_sc_hd__o22ai_4 _40593_ (.A1(_18108_),
    .A2(_18148_),
    .B1(_18213_),
    .B2(_18214_),
    .Y(_18215_));
 sky130_fd_sc_hd__a21o_1 _40594_ (.A1(_18201_),
    .A2(_18204_),
    .B1(_18212_),
    .X(_18216_));
 sky130_fd_sc_hd__nand3_4 _40595_ (.A(_18201_),
    .B(_18212_),
    .C(_18204_),
    .Y(_18217_));
 sky130_fd_sc_hd__nor2_2 _40596_ (.A(_18108_),
    .B(_18148_),
    .Y(_18218_));
 sky130_fd_sc_hd__nand3_4 _40597_ (.A(_18216_),
    .B(_18217_),
    .C(_18218_),
    .Y(_18219_));
 sky130_fd_sc_hd__nand2_1 _40598_ (.A(_18047_),
    .B(_17806_),
    .Y(_18220_));
 sky130_fd_sc_hd__nand2_2 _40599_ (.A(_18220_),
    .B(_18048_),
    .Y(_18221_));
 sky130_fd_sc_hd__nor2_2 _40600_ (.A(_17353_),
    .B(_18221_),
    .Y(_18222_));
 sky130_fd_sc_hd__and2_1 _40601_ (.A(_18221_),
    .B(_17353_),
    .X(_18223_));
 sky130_fd_sc_hd__nor2_2 _40602_ (.A(_18222_),
    .B(_18223_),
    .Y(_18224_));
 sky130_fd_sc_hd__a21oi_1 _40603_ (.A1(_18215_),
    .A2(_18219_),
    .B1(_18224_),
    .Y(_18225_));
 sky130_fd_sc_hd__nor2_2 _40604_ (.A(_16515_),
    .B(_18221_),
    .Y(_18226_));
 sky130_fd_sc_hd__nand2_1 _40605_ (.A(_18221_),
    .B(_17789_),
    .Y(_18227_));
 sky130_vsdinv _40606_ (.A(_18227_),
    .Y(_18228_));
 sky130_fd_sc_hd__o211a_1 _40607_ (.A1(_18226_),
    .A2(_18228_),
    .B1(_18219_),
    .C1(_18215_),
    .X(_18229_));
 sky130_fd_sc_hd__nand2_2 _40608_ (.A(_18134_),
    .B(_18119_),
    .Y(_18230_));
 sky130_fd_sc_hd__o21bai_1 _40609_ (.A1(_18225_),
    .A2(_18229_),
    .B1_N(_18230_),
    .Y(_18231_));
 sky130_fd_sc_hd__o2bb2ai_2 _40610_ (.A1_N(_18219_),
    .A2_N(_18215_),
    .B1(_18223_),
    .B2(_18222_),
    .Y(_18232_));
 sky130_fd_sc_hd__nand3_4 _40611_ (.A(_18215_),
    .B(_18219_),
    .C(_18224_),
    .Y(_18233_));
 sky130_fd_sc_hd__nand3_1 _40612_ (.A(_18232_),
    .B(_18233_),
    .C(_18230_),
    .Y(_18234_));
 sky130_fd_sc_hd__a21oi_1 _40613_ (.A1(_18231_),
    .A2(_18234_),
    .B1(_18125_),
    .Y(_18235_));
 sky130_vsdinv _40614_ (.A(_18125_),
    .Y(_18236_));
 sky130_fd_sc_hd__a21oi_4 _40615_ (.A1(_18232_),
    .A2(_18233_),
    .B1(_18230_),
    .Y(_18237_));
 sky130_fd_sc_hd__and3_2 _40616_ (.A(_18232_),
    .B(_18233_),
    .C(_18230_),
    .X(_18238_));
 sky130_fd_sc_hd__nor3_4 _40617_ (.A(_18236_),
    .B(_18237_),
    .C(_18238_),
    .Y(_18239_));
 sky130_fd_sc_hd__o21ai_2 _40618_ (.A1(_18139_),
    .A2(_18132_),
    .B1(_18138_),
    .Y(_18240_));
 sky130_fd_sc_hd__o21bai_2 _40619_ (.A1(_18235_),
    .A2(_18239_),
    .B1_N(_18240_),
    .Y(_18241_));
 sky130_fd_sc_hd__nor2_4 _40620_ (.A(_18236_),
    .B(_18237_),
    .Y(_18242_));
 sky130_fd_sc_hd__nand2_1 _40621_ (.A(_18242_),
    .B(_18234_),
    .Y(_18243_));
 sky130_fd_sc_hd__o21ai_2 _40622_ (.A1(_18237_),
    .A2(_18238_),
    .B1(_18236_),
    .Y(_18244_));
 sky130_fd_sc_hd__nand3_4 _40623_ (.A(_18243_),
    .B(_18240_),
    .C(_18244_),
    .Y(_18245_));
 sky130_fd_sc_hd__a21boi_4 _40624_ (.A1(_18143_),
    .A2(_18038_),
    .B1_N(_18144_),
    .Y(_18246_));
 sky130_fd_sc_hd__nor3_4 _40625_ (.A(_18139_),
    .B(_18132_),
    .C(_18135_),
    .Y(_18247_));
 sky130_fd_sc_hd__o22ai_1 _40626_ (.A1(_17789_),
    .A2(_18022_),
    .B1(_18132_),
    .B2(_18135_),
    .Y(_18248_));
 sky130_fd_sc_hd__nand2_1 _40627_ (.A(_18248_),
    .B(_18142_),
    .Y(_18249_));
 sky130_fd_sc_hd__o2111ai_4 _40628_ (.A1(_18247_),
    .A2(_18249_),
    .B1(_18035_),
    .C1(_18038_),
    .D1(_18144_),
    .Y(_18250_));
 sky130_fd_sc_hd__a21oi_4 _40629_ (.A1(_18041_),
    .A2(_18044_),
    .B1(_18250_),
    .Y(_18251_));
 sky130_fd_sc_hd__a211oi_4 _40630_ (.A1(_18241_),
    .A2(_18245_),
    .B1(_18246_),
    .C1(_18251_),
    .Y(_18252_));
 sky130_fd_sc_hd__nand2_1 _40631_ (.A(_18241_),
    .B(_18245_),
    .Y(_18253_));
 sky130_fd_sc_hd__o21bai_2 _40632_ (.A1(_18246_),
    .A2(_18251_),
    .B1_N(_18253_),
    .Y(_18254_));
 sky130_fd_sc_hd__nor2b_4 _40633_ (.A(_18252_),
    .B_N(_18254_),
    .Y(_02681_));
 sky130_fd_sc_hd__mux2_4 _40634_ (.A0(_16143_),
    .A1(_16142_),
    .S(_13989_),
    .X(_18255_));
 sky130_fd_sc_hd__xnor2_4 _40635_ (.A(_18255_),
    .B(_18173_),
    .Y(_18256_));
 sky130_fd_sc_hd__o21ai_4 _40636_ (.A1(_17436_),
    .A2(_18182_),
    .B1(_17434_),
    .Y(_18257_));
 sky130_fd_sc_hd__xor2_4 _40637_ (.A(_18066_),
    .B(_18257_),
    .X(_18258_));
 sky130_fd_sc_hd__xor2_4 _40638_ (.A(_18153_),
    .B(_18258_),
    .X(_18259_));
 sky130_fd_sc_hd__xor2_4 _40639_ (.A(_18256_),
    .B(_18259_),
    .X(_18260_));
 sky130_fd_sc_hd__nor3_4 _40640_ (.A(_18238_),
    .B(_18260_),
    .C(_18242_),
    .Y(_18261_));
 sky130_fd_sc_hd__o21a_1 _40641_ (.A1(_18238_),
    .A2(_18242_),
    .B1(_18260_),
    .X(_18262_));
 sky130_fd_sc_hd__nand2_2 _40642_ (.A(_18171_),
    .B(_18169_),
    .Y(_18263_));
 sky130_fd_sc_hd__nand2_2 _40643_ (.A(_18186_),
    .B(_18180_),
    .Y(_18264_));
 sky130_fd_sc_hd__xor2_4 _40644_ (.A(_18263_),
    .B(_18264_),
    .X(_18265_));
 sky130_fd_sc_hd__a21o_1 _40645_ (.A1(_18217_),
    .A2(_18204_),
    .B1(_18265_),
    .X(_18266_));
 sky130_fd_sc_hd__nand3_4 _40646_ (.A(_18217_),
    .B(_18204_),
    .C(_18265_),
    .Y(_18267_));
 sky130_fd_sc_hd__nand2_2 _40647_ (.A(_18179_),
    .B(_18165_),
    .Y(_18268_));
 sky130_fd_sc_hd__a21bo_1 _40648_ (.A1(_18190_),
    .A2(_18196_),
    .B1_N(_18187_),
    .X(_18269_));
 sky130_fd_sc_hd__xnor2_2 _40649_ (.A(_18268_),
    .B(_18269_),
    .Y(_18270_));
 sky130_fd_sc_hd__a21o_1 _40650_ (.A1(_18266_),
    .A2(_18267_),
    .B1(_18270_),
    .X(_18271_));
 sky130_fd_sc_hd__nand3_4 _40651_ (.A(_18266_),
    .B(_18270_),
    .C(_18267_),
    .Y(_18272_));
 sky130_fd_sc_hd__or2_1 _40652_ (.A(_17172_),
    .B(_18192_),
    .X(_18273_));
 sky130_fd_sc_hd__a21o_1 _40653_ (.A1(_18192_),
    .A2(_17162_),
    .B1(_16048_),
    .X(_18274_));
 sky130_fd_sc_hd__nor2_4 _40654_ (.A(_18154_),
    .B(_18156_),
    .Y(_18275_));
 sky130_fd_sc_hd__nand2_2 _40655_ (.A(_17245_),
    .B(_11294_),
    .Y(_18276_));
 sky130_fd_sc_hd__o21ai_4 _40656_ (.A1(_18152_),
    .A2(_18162_),
    .B1(_18161_),
    .Y(_18277_));
 sky130_fd_sc_hd__xor2_4 _40657_ (.A(_18276_),
    .B(_18277_),
    .X(_18278_));
 sky130_fd_sc_hd__xor2_4 _40658_ (.A(_18275_),
    .B(_18278_),
    .X(_18279_));
 sky130_fd_sc_hd__a21oi_2 _40659_ (.A1(_18273_),
    .A2(_18274_),
    .B1(_18279_),
    .Y(_18280_));
 sky130_fd_sc_hd__and3_1 _40660_ (.A(_18273_),
    .B(_18279_),
    .C(_18274_),
    .X(_18281_));
 sky130_fd_sc_hd__nor2_4 _40661_ (.A(_18280_),
    .B(_18281_),
    .Y(_18282_));
 sky130_fd_sc_hd__a21o_1 _40662_ (.A1(_18271_),
    .A2(_18272_),
    .B1(_18282_),
    .X(_18283_));
 sky130_fd_sc_hd__nand3_4 _40663_ (.A(_18271_),
    .B(_18282_),
    .C(_18272_),
    .Y(_18284_));
 sky130_fd_sc_hd__nand2_1 _40664_ (.A(_18283_),
    .B(_18284_),
    .Y(_18285_));
 sky130_fd_sc_hd__o21ai_1 _40665_ (.A1(_17891_),
    .A2(_18209_),
    .B1(_18208_),
    .Y(_18286_));
 sky130_fd_sc_hd__xnor2_1 _40666_ (.A(_18226_),
    .B(_18286_),
    .Y(_18287_));
 sky130_fd_sc_hd__nand3b_4 _40667_ (.A_N(_18287_),
    .B(_18233_),
    .C(_18219_),
    .Y(_18288_));
 sky130_fd_sc_hd__a21bo_1 _40668_ (.A1(_18233_),
    .A2(_18219_),
    .B1_N(_18287_),
    .X(_18289_));
 sky130_fd_sc_hd__nand3_4 _40669_ (.A(_18285_),
    .B(_18288_),
    .C(_18289_),
    .Y(_18290_));
 sky130_fd_sc_hd__nand2_1 _40670_ (.A(_18289_),
    .B(_18288_),
    .Y(_18291_));
 sky130_fd_sc_hd__nand3_4 _40671_ (.A(_18291_),
    .B(_18283_),
    .C(_18284_),
    .Y(_18292_));
 sky130_fd_sc_hd__nor2_8 _40672_ (.A(net465),
    .B(_16353_),
    .Y(_18293_));
 sky130_fd_sc_hd__nand3_2 _40673_ (.A(_18290_),
    .B(_18292_),
    .C(_18293_),
    .Y(_18294_));
 sky130_fd_sc_hd__a21o_1 _40674_ (.A1(_18290_),
    .A2(_18292_),
    .B1(_18293_),
    .X(_18295_));
 sky130_fd_sc_hd__o211a_1 _40675_ (.A1(_18261_),
    .A2(_18262_),
    .B1(_18294_),
    .C1(_18295_),
    .X(_18296_));
 sky130_fd_sc_hd__a21oi_1 _40676_ (.A1(_18290_),
    .A2(_18292_),
    .B1(_18293_),
    .Y(_18297_));
 sky130_fd_sc_hd__and3_1 _40677_ (.A(_18290_),
    .B(_18292_),
    .C(_18293_),
    .X(_18298_));
 sky130_fd_sc_hd__nor2_1 _40678_ (.A(_18261_),
    .B(_18262_),
    .Y(_18299_));
 sky130_fd_sc_hd__o21a_1 _40679_ (.A1(_18297_),
    .A2(_18298_),
    .B1(_18299_),
    .X(_18300_));
 sky130_fd_sc_hd__o2bb2ai_1 _40680_ (.A1_N(_18245_),
    .A2_N(_18254_),
    .B1(_18296_),
    .B2(_18300_),
    .Y(_18301_));
 sky130_fd_sc_hd__o22ai_1 _40681_ (.A1(_18262_),
    .A2(_18261_),
    .B1(_18297_),
    .B2(_18298_),
    .Y(_18302_));
 sky130_fd_sc_hd__nand3_1 _40682_ (.A(_18299_),
    .B(_18295_),
    .C(_18294_),
    .Y(_18303_));
 sky130_fd_sc_hd__nand2_1 _40683_ (.A(_18302_),
    .B(_18303_),
    .Y(_18304_));
 sky130_fd_sc_hd__nand3_1 _40684_ (.A(_18304_),
    .B(_18245_),
    .C(_18254_),
    .Y(_18305_));
 sky130_fd_sc_hd__nand2_2 _40685_ (.A(_18301_),
    .B(_18305_),
    .Y(_02682_));
 sky130_fd_sc_hd__xnor2_1 _40686_ (.A(_05349_),
    .B(_05196_),
    .Y(_02628_));
 sky130_fd_sc_hd__nor2_1 _40687_ (.A(_20119_),
    .B(_04847_),
    .Y(_00050_));
 sky130_fd_sc_hd__and2_1 _40688_ (.A(_02318_),
    .B(_00066_),
    .X(_00067_));
 sky130_fd_sc_hd__and2_1 _40689_ (.A(_02321_),
    .B(_00084_),
    .X(_00085_));
 sky130_fd_sc_hd__and2_1 _40690_ (.A(_02321_),
    .B(_00094_),
    .X(_00095_));
 sky130_fd_sc_hd__o21a_4 _40691_ (.A1(instr_sra),
    .A2(instr_srai),
    .B1(_18451_),
    .X(_00216_));
 sky130_fd_sc_hd__o21a_1 _40692_ (.A1(_18525_),
    .A2(_18535_),
    .B1(_00321_),
    .X(_18306_));
 sky130_fd_sc_hd__nand2_1 _40693_ (.A(_18306_),
    .B(_18496_),
    .Y(_18307_));
 sky130_fd_sc_hd__o211a_1 _40694_ (.A1(irq_active),
    .A2(_18306_),
    .B1(_18938_),
    .C1(_18307_),
    .X(_04072_));
 sky130_fd_sc_hd__conb_1 _40695_ (.LO(net134));
 sky130_fd_sc_hd__conb_1 _40696_ (.LO(net145));
 sky130_fd_sc_hd__conb_1 _40697_ (.LO(net167));
 sky130_fd_sc_hd__conb_1 _40698_ (.LO(net178));
 sky130_fd_sc_hd__conb_1 _40699_ (.LO(net371));
 sky130_fd_sc_hd__conb_1 _40700_ (.LO(net382));
 sky130_fd_sc_hd__conb_1 _40701_ (.LO(net393));
 sky130_fd_sc_hd__conb_1 _40702_ (.LO(net400));
 sky130_fd_sc_hd__conb_1 _40703_ (.LO(net401));
 sky130_fd_sc_hd__conb_1 _40704_ (.LO(net402));
 sky130_fd_sc_hd__conb_1 _40705_ (.LO(net403));
 sky130_fd_sc_hd__conb_1 _40706_ (.LO(net404));
 sky130_fd_sc_hd__conb_1 _40707_ (.LO(net405));
 sky130_fd_sc_hd__conb_1 _40708_ (.LO(net406));
 sky130_fd_sc_hd__conb_1 _40709_ (.LO(net372));
 sky130_fd_sc_hd__conb_1 _40710_ (.LO(net373));
 sky130_fd_sc_hd__conb_1 _40711_ (.LO(net374));
 sky130_fd_sc_hd__conb_1 _40712_ (.LO(net375));
 sky130_fd_sc_hd__conb_1 _40713_ (.LO(net376));
 sky130_fd_sc_hd__conb_1 _40714_ (.LO(net377));
 sky130_fd_sc_hd__conb_1 _40715_ (.LO(net378));
 sky130_fd_sc_hd__conb_1 _40716_ (.LO(net379));
 sky130_fd_sc_hd__conb_1 _40717_ (.LO(net380));
 sky130_fd_sc_hd__conb_1 _40718_ (.LO(net381));
 sky130_fd_sc_hd__conb_1 _40719_ (.LO(net383));
 sky130_fd_sc_hd__conb_1 _40720_ (.LO(net384));
 sky130_fd_sc_hd__conb_1 _40721_ (.LO(net385));
 sky130_fd_sc_hd__conb_1 _40722_ (.LO(net386));
 sky130_fd_sc_hd__conb_1 _40723_ (.LO(net387));
 sky130_fd_sc_hd__conb_1 _40724_ (.LO(net388));
 sky130_fd_sc_hd__conb_1 _40725_ (.LO(net389));
 sky130_fd_sc_hd__conb_1 _40726_ (.LO(net390));
 sky130_fd_sc_hd__conb_1 _40727_ (.LO(net391));
 sky130_fd_sc_hd__conb_1 _40728_ (.LO(net392));
 sky130_fd_sc_hd__conb_1 _40729_ (.LO(net394));
 sky130_fd_sc_hd__conb_1 _40730_ (.LO(net395));
 sky130_fd_sc_hd__conb_1 _40731_ (.LO(net396));
 sky130_fd_sc_hd__conb_1 _40732_ (.LO(net397));
 sky130_fd_sc_hd__conb_1 _40733_ (.LO(net398));
 sky130_fd_sc_hd__conb_1 _40734_ (.LO(net399));
 sky130_fd_sc_hd__conb_1 _40735_ (.LO(net407));
 sky130_fd_sc_hd__conb_1 _40736_ (.LO(_00313_));
 sky130_fd_sc_hd__buf_4 _40737_ (.A(net200),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 _40738_ (.A(net211),
    .X(net349));
 sky130_fd_sc_hd__buf_6 _40739_ (.A(net222),
    .X(net360));
 sky130_fd_sc_hd__buf_2 _40740_ (.A(net225),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 _40741_ (.A(net502),
    .X(net364));
 sky130_fd_sc_hd__buf_2 _40742_ (.A(net227),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 _40743_ (.A(net228),
    .X(net366));
 sky130_fd_sc_hd__buf_2 _40744_ (.A(net229),
    .X(net367));
 sky130_fd_sc_hd__mux2_8 _40745_ (.A0(decoder_trigger),
    .A1(_02410_),
    .S(_00309_),
    .X(_20894_));
 sky130_fd_sc_hd__mux2_1 _40746_ (.A0(\reg_out[2] ),
    .A1(\reg_next_pc[2] ),
    .S(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_8 _40747_ (.A0(_02184_),
    .A1(net328),
    .S(net462),
    .X(net189));
 sky130_fd_sc_hd__mux2_2 _40748_ (.A0(\reg_out[3] ),
    .A1(\reg_next_pc[3] ),
    .S(_02183_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_4 _40749_ (.A0(_02185_),
    .A1(net331),
    .S(net460),
    .X(net192));
 sky130_fd_sc_hd__mux2_1 _40750_ (.A0(\reg_out[4] ),
    .A1(\reg_next_pc[4] ),
    .S(_02183_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_8 _40751_ (.A0(_02186_),
    .A1(net332),
    .S(net462),
    .X(net193));
 sky130_fd_sc_hd__mux2_1 _40752_ (.A0(\reg_out[5] ),
    .A1(\reg_next_pc[5] ),
    .S(_02183_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_8 _40753_ (.A0(_02187_),
    .A1(net333),
    .S(net461),
    .X(net194));
 sky130_fd_sc_hd__mux2_4 _40754_ (.A0(\reg_out[6] ),
    .A1(\reg_next_pc[6] ),
    .S(_02183_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_4 _40755_ (.A0(_02188_),
    .A1(net334),
    .S(net460),
    .X(net195));
 sky130_fd_sc_hd__mux2_2 _40756_ (.A0(\reg_out[7] ),
    .A1(\reg_next_pc[7] ),
    .S(_02183_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_4 _40757_ (.A0(_02189_),
    .A1(net335),
    .S(net460),
    .X(net196));
 sky130_fd_sc_hd__mux2_2 _40758_ (.A0(\reg_out[8] ),
    .A1(\reg_next_pc[8] ),
    .S(_02183_),
    .X(_02190_));
 sky130_fd_sc_hd__mux2_4 _40759_ (.A0(_02190_),
    .A1(net336),
    .S(net460),
    .X(net197));
 sky130_fd_sc_hd__mux2_1 _40760_ (.A0(\reg_out[9] ),
    .A1(\reg_next_pc[9] ),
    .S(_02183_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_8 _40761_ (.A0(_02191_),
    .A1(net337),
    .S(net459),
    .X(net198));
 sky130_fd_sc_hd__mux2_1 _40762_ (.A0(\reg_out[10] ),
    .A1(\reg_next_pc[10] ),
    .S(_02183_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_8 _40763_ (.A0(_02192_),
    .A1(net307),
    .S(net461),
    .X(net168));
 sky130_fd_sc_hd__mux2_1 _40764_ (.A0(\reg_out[11] ),
    .A1(\reg_next_pc[11] ),
    .S(_02183_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_8 _40765_ (.A0(_02193_),
    .A1(net308),
    .S(net460),
    .X(net169));
 sky130_fd_sc_hd__mux2_1 _40766_ (.A0(\reg_out[12] ),
    .A1(\reg_next_pc[12] ),
    .S(_02183_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_8 _40767_ (.A0(_02194_),
    .A1(net309),
    .S(net461),
    .X(net170));
 sky130_fd_sc_hd__mux2_4 _40768_ (.A0(\reg_out[13] ),
    .A1(\reg_next_pc[13] ),
    .S(_02183_),
    .X(_02195_));
 sky130_fd_sc_hd__mux2_8 _40769_ (.A0(_02195_),
    .A1(net310),
    .S(net460),
    .X(net171));
 sky130_fd_sc_hd__mux2_1 _40770_ (.A0(\reg_out[14] ),
    .A1(\reg_next_pc[14] ),
    .S(_02183_),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_8 _40771_ (.A0(_02196_),
    .A1(net311),
    .S(net459),
    .X(net172));
 sky130_fd_sc_hd__mux2_1 _40772_ (.A0(\reg_out[15] ),
    .A1(\reg_next_pc[15] ),
    .S(_02183_),
    .X(_02197_));
 sky130_fd_sc_hd__mux2_2 _40773_ (.A0(_02197_),
    .A1(net312),
    .S(net461),
    .X(net173));
 sky130_fd_sc_hd__mux2_1 _40774_ (.A0(\reg_out[16] ),
    .A1(\reg_next_pc[16] ),
    .S(_02183_),
    .X(_02198_));
 sky130_fd_sc_hd__mux2_8 _40775_ (.A0(_02198_),
    .A1(net313),
    .S(net459),
    .X(net174));
 sky130_fd_sc_hd__mux2_1 _40776_ (.A0(\reg_out[17] ),
    .A1(\reg_next_pc[17] ),
    .S(_02183_),
    .X(_02199_));
 sky130_fd_sc_hd__mux2_8 _40777_ (.A0(_02199_),
    .A1(net314),
    .S(net459),
    .X(net175));
 sky130_fd_sc_hd__mux2_1 _40778_ (.A0(\reg_out[18] ),
    .A1(\reg_next_pc[18] ),
    .S(_02183_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_8 _40779_ (.A0(_02200_),
    .A1(net315),
    .S(net459),
    .X(net176));
 sky130_fd_sc_hd__mux2_1 _40780_ (.A0(\reg_out[19] ),
    .A1(\reg_next_pc[19] ),
    .S(_02183_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_8 _40781_ (.A0(_02201_),
    .A1(net316),
    .S(net459),
    .X(net177));
 sky130_fd_sc_hd__mux2_4 _40782_ (.A0(\reg_out[20] ),
    .A1(\reg_next_pc[20] ),
    .S(_02183_),
    .X(_02202_));
 sky130_fd_sc_hd__mux2_4 _40783_ (.A0(_02202_),
    .A1(net318),
    .S(net460),
    .X(net179));
 sky130_fd_sc_hd__mux2_1 _40784_ (.A0(\reg_out[21] ),
    .A1(\reg_next_pc[21] ),
    .S(_02183_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_8 _40785_ (.A0(_02203_),
    .A1(net319),
    .S(net459),
    .X(net180));
 sky130_fd_sc_hd__mux2_1 _40786_ (.A0(\reg_out[22] ),
    .A1(\reg_next_pc[22] ),
    .S(_02183_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_8 _40787_ (.A0(_02204_),
    .A1(net320),
    .S(net459),
    .X(net181));
 sky130_fd_sc_hd__mux2_2 _40788_ (.A0(\reg_out[23] ),
    .A1(\reg_next_pc[23] ),
    .S(_02183_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_8 _40789_ (.A0(_02205_),
    .A1(net321),
    .S(net461),
    .X(net182));
 sky130_fd_sc_hd__mux2_2 _40790_ (.A0(\reg_out[24] ),
    .A1(\reg_next_pc[24] ),
    .S(_02183_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_8 _40791_ (.A0(_02206_),
    .A1(net322),
    .S(net461),
    .X(net183));
 sky130_fd_sc_hd__mux2_4 _40792_ (.A0(\reg_out[25] ),
    .A1(\reg_next_pc[25] ),
    .S(_02183_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_2 _40793_ (.A0(_02207_),
    .A1(net323),
    .S(net460),
    .X(net184));
 sky130_fd_sc_hd__mux2_1 _40794_ (.A0(\reg_out[26] ),
    .A1(\reg_next_pc[26] ),
    .S(_02183_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_8 _40795_ (.A0(_02208_),
    .A1(net324),
    .S(net462),
    .X(net185));
 sky130_fd_sc_hd__mux2_1 _40796_ (.A0(\reg_out[27] ),
    .A1(\reg_next_pc[27] ),
    .S(_02183_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_4 _40797_ (.A0(_02209_),
    .A1(net325),
    .S(net462),
    .X(net186));
 sky130_fd_sc_hd__mux2_2 _40798_ (.A0(\reg_out[28] ),
    .A1(\reg_next_pc[28] ),
    .S(_02183_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_8 _40799_ (.A0(_02210_),
    .A1(net326),
    .S(net461),
    .X(net187));
 sky130_fd_sc_hd__mux2_1 _40800_ (.A0(\reg_out[29] ),
    .A1(\reg_next_pc[29] ),
    .S(_02183_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_8 _40801_ (.A0(_02211_),
    .A1(net327),
    .S(net462),
    .X(net188));
 sky130_fd_sc_hd__mux2_1 _40802_ (.A0(\reg_out[30] ),
    .A1(\reg_next_pc[30] ),
    .S(_02183_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_8 _40803_ (.A0(_02212_),
    .A1(net329),
    .S(net462),
    .X(net190));
 sky130_fd_sc_hd__mux2_4 _40804_ (.A0(\reg_out[31] ),
    .A1(\reg_next_pc[31] ),
    .S(_02183_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_2 _40805_ (.A0(_02213_),
    .A1(net330),
    .S(net460),
    .X(net191));
 sky130_fd_sc_hd__mux2_8 _40806_ (.A0(_02167_),
    .A1(net368),
    .S(net432),
    .X(net230));
 sky130_fd_sc_hd__mux2_8 _40807_ (.A0(_02168_),
    .A1(net369),
    .S(net433),
    .X(net231));
 sky130_fd_sc_hd__mux2_8 _40808_ (.A0(_02169_),
    .A1(net339),
    .S(net433),
    .X(net201));
 sky130_fd_sc_hd__mux2_8 _40809_ (.A0(_02170_),
    .A1(net340),
    .S(net433),
    .X(net202));
 sky130_fd_sc_hd__mux2_8 _40810_ (.A0(_02171_),
    .A1(net341),
    .S(net433),
    .X(net203));
 sky130_fd_sc_hd__mux2_4 _40811_ (.A0(_02172_),
    .A1(net342),
    .S(_01683_),
    .X(net204));
 sky130_fd_sc_hd__mux2_8 _40812_ (.A0(_02173_),
    .A1(net343),
    .S(net433),
    .X(net205));
 sky130_fd_sc_hd__mux2_8 _40813_ (.A0(_02174_),
    .A1(net344),
    .S(net432),
    .X(net206));
 sky130_fd_sc_hd__mux2_8 _40814_ (.A0(_02175_),
    .A1(net345),
    .S(net432),
    .X(net207));
 sky130_fd_sc_hd__mux2_8 _40815_ (.A0(_02176_),
    .A1(net346),
    .S(net434),
    .X(net208));
 sky130_fd_sc_hd__mux2_8 _40816_ (.A0(_02177_),
    .A1(net347),
    .S(_01683_),
    .X(net209));
 sky130_fd_sc_hd__mux2_8 _40817_ (.A0(_02178_),
    .A1(net348),
    .S(net434),
    .X(net210));
 sky130_fd_sc_hd__mux2_8 _40818_ (.A0(_02179_),
    .A1(net350),
    .S(net434),
    .X(net212));
 sky130_fd_sc_hd__mux2_8 _40819_ (.A0(_02180_),
    .A1(net351),
    .S(net434),
    .X(net213));
 sky130_fd_sc_hd__mux2_8 _40820_ (.A0(_02181_),
    .A1(net352),
    .S(net434),
    .X(net214));
 sky130_fd_sc_hd__mux2_8 _40821_ (.A0(_02182_),
    .A1(net353),
    .S(net434),
    .X(net215));
 sky130_fd_sc_hd__mux2_8 _40822_ (.A0(_02167_),
    .A1(net354),
    .S(net432),
    .X(net216));
 sky130_fd_sc_hd__mux2_8 _40823_ (.A0(_02168_),
    .A1(net355),
    .S(net433),
    .X(net217));
 sky130_fd_sc_hd__mux2_8 _40824_ (.A0(_02169_),
    .A1(net356),
    .S(net433),
    .X(net218));
 sky130_fd_sc_hd__mux2_8 _40825_ (.A0(_02170_),
    .A1(net357),
    .S(_01683_),
    .X(net219));
 sky130_fd_sc_hd__mux2_8 _40826_ (.A0(_02171_),
    .A1(net358),
    .S(net432),
    .X(net220));
 sky130_fd_sc_hd__mux2_8 _40827_ (.A0(_02172_),
    .A1(net359),
    .S(_01683_),
    .X(net221));
 sky130_fd_sc_hd__mux2_8 _40828_ (.A0(_02173_),
    .A1(net361),
    .S(net433),
    .X(net223));
 sky130_fd_sc_hd__mux2_8 _40829_ (.A0(_02174_),
    .A1(net362),
    .S(net432),
    .X(net224));
 sky130_fd_sc_hd__mux2_1 _40830_ (.A0(\mem_rdata_q[7] ),
    .A1(net62),
    .S(net479),
    .X(\mem_rdata_latched[7] ));
 sky130_fd_sc_hd__mux2_1 _40831_ (.A0(\mem_rdata_q[8] ),
    .A1(net63),
    .S(net479),
    .X(\mem_rdata_latched[8] ));
 sky130_fd_sc_hd__mux2_1 _40832_ (.A0(\mem_rdata_q[9] ),
    .A1(net64),
    .S(net479),
    .X(\mem_rdata_latched[9] ));
 sky130_fd_sc_hd__mux2_1 _40833_ (.A0(\mem_rdata_q[10] ),
    .A1(net34),
    .S(net479),
    .X(\mem_rdata_latched[10] ));
 sky130_fd_sc_hd__mux2_1 _40834_ (.A0(\mem_rdata_q[11] ),
    .A1(net35),
    .S(net479),
    .X(\mem_rdata_latched[11] ));
 sky130_fd_sc_hd__mux2_2 _40835_ (.A0(\mem_rdata_q[12] ),
    .A1(net517),
    .S(net479),
    .X(\mem_rdata_latched[12] ));
 sky130_fd_sc_hd__mux2_2 _40836_ (.A0(\mem_rdata_q[13] ),
    .A1(net37),
    .S(net479),
    .X(\mem_rdata_latched[13] ));
 sky130_fd_sc_hd__mux2_2 _40837_ (.A0(\mem_rdata_q[14] ),
    .A1(net38),
    .S(net479),
    .X(\mem_rdata_latched[14] ));
 sky130_fd_sc_hd__mux2_1 _40838_ (.A0(\mem_rdata_q[15] ),
    .A1(net516),
    .S(net479),
    .X(\mem_rdata_latched[15] ));
 sky130_fd_sc_hd__mux2_1 _40839_ (.A0(\mem_rdata_q[16] ),
    .A1(net40),
    .S(net479),
    .X(\mem_rdata_latched[16] ));
 sky130_fd_sc_hd__mux2_1 _40840_ (.A0(\mem_rdata_q[17] ),
    .A1(net41),
    .S(net479),
    .X(\mem_rdata_latched[17] ));
 sky130_fd_sc_hd__mux2_1 _40841_ (.A0(\mem_rdata_q[18] ),
    .A1(net42),
    .S(net479),
    .X(\mem_rdata_latched[18] ));
 sky130_fd_sc_hd__mux2_1 _40842_ (.A0(\mem_rdata_q[19] ),
    .A1(net515),
    .S(net479),
    .X(\mem_rdata_latched[19] ));
 sky130_fd_sc_hd__mux2_1 _40843_ (.A0(\mem_rdata_q[20] ),
    .A1(net514),
    .S(net479),
    .X(\mem_rdata_latched[20] ));
 sky130_fd_sc_hd__mux2_1 _40844_ (.A0(\mem_rdata_q[21] ),
    .A1(net46),
    .S(net479),
    .X(\mem_rdata_latched[21] ));
 sky130_fd_sc_hd__mux2_1 _40845_ (.A0(\mem_rdata_q[22] ),
    .A1(net47),
    .S(net479),
    .X(\mem_rdata_latched[22] ));
 sky130_fd_sc_hd__mux2_1 _40846_ (.A0(\mem_rdata_q[23] ),
    .A1(net48),
    .S(net479),
    .X(\mem_rdata_latched[23] ));
 sky130_fd_sc_hd__mux2_1 _40847_ (.A0(\mem_rdata_q[24] ),
    .A1(net49),
    .S(net479),
    .X(\mem_rdata_latched[24] ));
 sky130_fd_sc_hd__mux2_1 _40848_ (.A0(\mem_rdata_q[25] ),
    .A1(net50),
    .S(net479),
    .X(\mem_rdata_latched[25] ));
 sky130_fd_sc_hd__mux2_1 _40849_ (.A0(\mem_rdata_q[26] ),
    .A1(net51),
    .S(net479),
    .X(\mem_rdata_latched[26] ));
 sky130_fd_sc_hd__mux2_1 _40850_ (.A0(\mem_rdata_q[27] ),
    .A1(net52),
    .S(mem_xfer),
    .X(\mem_rdata_latched[27] ));
 sky130_fd_sc_hd__mux2_2 _40851_ (.A0(\mem_rdata_q[28] ),
    .A1(net53),
    .S(net479),
    .X(\mem_rdata_latched[28] ));
 sky130_fd_sc_hd__mux2_1 _40852_ (.A0(\mem_rdata_q[29] ),
    .A1(net54),
    .S(net479),
    .X(\mem_rdata_latched[29] ));
 sky130_fd_sc_hd__mux2_1 _40853_ (.A0(\mem_rdata_q[30] ),
    .A1(net513),
    .S(net479),
    .X(\mem_rdata_latched[30] ));
 sky130_fd_sc_hd__mux2_1 _40854_ (.A0(\mem_rdata_q[31] ),
    .A1(net57),
    .S(net479),
    .X(\mem_rdata_latched[31] ));
 sky130_fd_sc_hd__mux2_1 _40855_ (.A0(_02134_),
    .A1(\alu_add_sub[0] ),
    .S(_02133_),
    .X(\alu_out[0] ));
 sky130_fd_sc_hd__mux2_1 _40856_ (.A0(_02135_),
    .A1(\alu_add_sub[1] ),
    .S(_02133_),
    .X(\alu_out[1] ));
 sky130_fd_sc_hd__mux2_1 _40857_ (.A0(_02136_),
    .A1(\alu_add_sub[2] ),
    .S(_02133_),
    .X(\alu_out[2] ));
 sky130_fd_sc_hd__mux2_1 _40858_ (.A0(_02137_),
    .A1(\alu_add_sub[3] ),
    .S(_02133_),
    .X(\alu_out[3] ));
 sky130_fd_sc_hd__mux2_1 _40859_ (.A0(_02138_),
    .A1(\alu_add_sub[4] ),
    .S(_02133_),
    .X(\alu_out[4] ));
 sky130_fd_sc_hd__mux2_1 _40860_ (.A0(_02139_),
    .A1(\alu_add_sub[5] ),
    .S(_02133_),
    .X(\alu_out[5] ));
 sky130_fd_sc_hd__mux2_1 _40861_ (.A0(_02140_),
    .A1(\alu_add_sub[6] ),
    .S(_02133_),
    .X(\alu_out[6] ));
 sky130_fd_sc_hd__mux2_1 _40862_ (.A0(_02141_),
    .A1(\alu_add_sub[7] ),
    .S(_02133_),
    .X(\alu_out[7] ));
 sky130_fd_sc_hd__mux2_1 _40863_ (.A0(_02142_),
    .A1(\alu_add_sub[8] ),
    .S(_02133_),
    .X(\alu_out[8] ));
 sky130_fd_sc_hd__mux2_1 _40864_ (.A0(_02143_),
    .A1(\alu_add_sub[9] ),
    .S(_02133_),
    .X(\alu_out[9] ));
 sky130_fd_sc_hd__mux2_1 _40865_ (.A0(_02144_),
    .A1(\alu_add_sub[10] ),
    .S(_02133_),
    .X(\alu_out[10] ));
 sky130_fd_sc_hd__mux2_1 _40866_ (.A0(_02145_),
    .A1(\alu_add_sub[11] ),
    .S(_02133_),
    .X(\alu_out[11] ));
 sky130_fd_sc_hd__mux2_1 _40867_ (.A0(_02146_),
    .A1(\alu_add_sub[12] ),
    .S(_02133_),
    .X(\alu_out[12] ));
 sky130_fd_sc_hd__mux2_1 _40868_ (.A0(_02147_),
    .A1(\alu_add_sub[13] ),
    .S(_02133_),
    .X(\alu_out[13] ));
 sky130_fd_sc_hd__mux2_1 _40869_ (.A0(_02148_),
    .A1(\alu_add_sub[14] ),
    .S(_02133_),
    .X(\alu_out[14] ));
 sky130_fd_sc_hd__mux2_1 _40870_ (.A0(_02149_),
    .A1(\alu_add_sub[15] ),
    .S(_02133_),
    .X(\alu_out[15] ));
 sky130_fd_sc_hd__mux2_1 _40871_ (.A0(_02150_),
    .A1(\alu_add_sub[16] ),
    .S(_02133_),
    .X(\alu_out[16] ));
 sky130_fd_sc_hd__mux2_1 _40872_ (.A0(_02151_),
    .A1(\alu_add_sub[17] ),
    .S(_02133_),
    .X(\alu_out[17] ));
 sky130_fd_sc_hd__mux2_1 _40873_ (.A0(_02152_),
    .A1(\alu_add_sub[18] ),
    .S(_02133_),
    .X(\alu_out[18] ));
 sky130_fd_sc_hd__mux2_1 _40874_ (.A0(_02153_),
    .A1(\alu_add_sub[19] ),
    .S(_02133_),
    .X(\alu_out[19] ));
 sky130_fd_sc_hd__mux2_1 _40875_ (.A0(_02154_),
    .A1(\alu_add_sub[20] ),
    .S(_02133_),
    .X(\alu_out[20] ));
 sky130_fd_sc_hd__mux2_1 _40876_ (.A0(_02155_),
    .A1(\alu_add_sub[21] ),
    .S(_02133_),
    .X(\alu_out[21] ));
 sky130_fd_sc_hd__mux2_1 _40877_ (.A0(_02156_),
    .A1(\alu_add_sub[22] ),
    .S(_02133_),
    .X(\alu_out[22] ));
 sky130_fd_sc_hd__mux2_2 _40878_ (.A0(_02157_),
    .A1(\alu_add_sub[23] ),
    .S(_02133_),
    .X(\alu_out[23] ));
 sky130_fd_sc_hd__mux2_2 _40879_ (.A0(_02158_),
    .A1(\alu_add_sub[24] ),
    .S(_02133_),
    .X(\alu_out[24] ));
 sky130_fd_sc_hd__mux2_2 _40880_ (.A0(_02159_),
    .A1(\alu_add_sub[25] ),
    .S(_02133_),
    .X(\alu_out[25] ));
 sky130_fd_sc_hd__mux2_1 _40881_ (.A0(_02160_),
    .A1(\alu_add_sub[26] ),
    .S(_02133_),
    .X(\alu_out[26] ));
 sky130_fd_sc_hd__mux2_1 _40882_ (.A0(_02161_),
    .A1(\alu_add_sub[27] ),
    .S(_02133_),
    .X(\alu_out[27] ));
 sky130_fd_sc_hd__mux2_1 _40883_ (.A0(_02162_),
    .A1(\alu_add_sub[28] ),
    .S(_02133_),
    .X(\alu_out[28] ));
 sky130_fd_sc_hd__mux2_1 _40884_ (.A0(_02163_),
    .A1(\alu_add_sub[29] ),
    .S(_02133_),
    .X(\alu_out[29] ));
 sky130_fd_sc_hd__mux2_1 _40885_ (.A0(_02164_),
    .A1(\alu_add_sub[30] ),
    .S(_02133_),
    .X(\alu_out[30] ));
 sky130_fd_sc_hd__mux2_1 _40886_ (.A0(_02165_),
    .A1(\alu_add_sub[31] ),
    .S(_02133_),
    .X(\alu_out[31] ));
 sky130_fd_sc_hd__mux2_4 _40887_ (.A0(_02071_),
    .A1(\reg_next_pc[0] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[0] ));
 sky130_fd_sc_hd__mux2_4 _40888_ (.A0(_02072_),
    .A1(\reg_pc[1] ),
    .S(_02069_),
    .X(\cpuregs_wrdata[1] ));
 sky130_fd_sc_hd__mux2_4 _40889_ (.A0(_02074_),
    .A1(_02073_),
    .S(_02069_),
    .X(\cpuregs_wrdata[2] ));
 sky130_fd_sc_hd__mux2_4 _40890_ (.A0(_02076_),
    .A1(_02075_),
    .S(_02069_),
    .X(\cpuregs_wrdata[3] ));
 sky130_fd_sc_hd__mux2_4 _40891_ (.A0(_02078_),
    .A1(_02077_),
    .S(_02069_),
    .X(\cpuregs_wrdata[4] ));
 sky130_fd_sc_hd__mux2_4 _40892_ (.A0(_02080_),
    .A1(_02079_),
    .S(_02069_),
    .X(\cpuregs_wrdata[5] ));
 sky130_fd_sc_hd__mux2_4 _40893_ (.A0(_02082_),
    .A1(_02081_),
    .S(net429),
    .X(\cpuregs_wrdata[6] ));
 sky130_fd_sc_hd__mux2_4 _40894_ (.A0(_02084_),
    .A1(_02083_),
    .S(net429),
    .X(\cpuregs_wrdata[7] ));
 sky130_fd_sc_hd__mux2_4 _40895_ (.A0(_02086_),
    .A1(_02085_),
    .S(net429),
    .X(\cpuregs_wrdata[8] ));
 sky130_fd_sc_hd__mux2_4 _40896_ (.A0(_02088_),
    .A1(_02087_),
    .S(net429),
    .X(\cpuregs_wrdata[9] ));
 sky130_fd_sc_hd__mux2_4 _40897_ (.A0(_02090_),
    .A1(_02089_),
    .S(net429),
    .X(\cpuregs_wrdata[10] ));
 sky130_fd_sc_hd__mux2_4 _40898_ (.A0(_02092_),
    .A1(_02091_),
    .S(net429),
    .X(\cpuregs_wrdata[11] ));
 sky130_fd_sc_hd__mux2_4 _40899_ (.A0(_02094_),
    .A1(_02093_),
    .S(net429),
    .X(\cpuregs_wrdata[12] ));
 sky130_fd_sc_hd__mux2_4 _40900_ (.A0(_02096_),
    .A1(_02095_),
    .S(net429),
    .X(\cpuregs_wrdata[13] ));
 sky130_fd_sc_hd__mux2_2 _40901_ (.A0(_02098_),
    .A1(_02097_),
    .S(net429),
    .X(\cpuregs_wrdata[14] ));
 sky130_fd_sc_hd__mux2_2 _40902_ (.A0(_02100_),
    .A1(_02099_),
    .S(net429),
    .X(\cpuregs_wrdata[15] ));
 sky130_fd_sc_hd__mux2_2 _40903_ (.A0(_02102_),
    .A1(_02101_),
    .S(net429),
    .X(\cpuregs_wrdata[16] ));
 sky130_fd_sc_hd__mux2_2 _40904_ (.A0(_02104_),
    .A1(_02103_),
    .S(net429),
    .X(\cpuregs_wrdata[17] ));
 sky130_fd_sc_hd__mux2_2 _40905_ (.A0(_02106_),
    .A1(_02105_),
    .S(net430),
    .X(\cpuregs_wrdata[18] ));
 sky130_fd_sc_hd__mux2_2 _40906_ (.A0(_02108_),
    .A1(_02107_),
    .S(net430),
    .X(\cpuregs_wrdata[19] ));
 sky130_fd_sc_hd__mux2_4 _40907_ (.A0(_02110_),
    .A1(_02109_),
    .S(net430),
    .X(\cpuregs_wrdata[20] ));
 sky130_fd_sc_hd__mux2_2 _40908_ (.A0(_02112_),
    .A1(_02111_),
    .S(net430),
    .X(\cpuregs_wrdata[21] ));
 sky130_fd_sc_hd__mux2_2 _40909_ (.A0(_02114_),
    .A1(_02113_),
    .S(net430),
    .X(\cpuregs_wrdata[22] ));
 sky130_fd_sc_hd__mux2_4 _40910_ (.A0(_02116_),
    .A1(_02115_),
    .S(net430),
    .X(\cpuregs_wrdata[23] ));
 sky130_fd_sc_hd__mux2_4 _40911_ (.A0(_02118_),
    .A1(_02117_),
    .S(net430),
    .X(\cpuregs_wrdata[24] ));
 sky130_fd_sc_hd__mux2_4 _40912_ (.A0(_02120_),
    .A1(_02119_),
    .S(net430),
    .X(\cpuregs_wrdata[25] ));
 sky130_fd_sc_hd__mux2_2 _40913_ (.A0(_02122_),
    .A1(_02121_),
    .S(_02069_),
    .X(\cpuregs_wrdata[26] ));
 sky130_fd_sc_hd__mux2_4 _40914_ (.A0(_02124_),
    .A1(_02123_),
    .S(_02069_),
    .X(\cpuregs_wrdata[27] ));
 sky130_fd_sc_hd__mux2_4 _40915_ (.A0(_02126_),
    .A1(_02125_),
    .S(_02069_),
    .X(\cpuregs_wrdata[28] ));
 sky130_fd_sc_hd__mux2_4 _40916_ (.A0(_02128_),
    .A1(_02127_),
    .S(_02069_),
    .X(\cpuregs_wrdata[29] ));
 sky130_fd_sc_hd__mux2_4 _40917_ (.A0(_02130_),
    .A1(_02129_),
    .S(_02069_),
    .X(\cpuregs_wrdata[30] ));
 sky130_fd_sc_hd__mux2_2 _40918_ (.A0(_02132_),
    .A1(_02131_),
    .S(_02069_),
    .X(\cpuregs_wrdata[31] ));
 sky130_fd_sc_hd__mux2_1 _40919_ (.A0(_02316_),
    .A1(_02317_),
    .S(_00307_),
    .X(_00004_));
 sky130_fd_sc_hd__mux2_1 _40920_ (.A0(_00347_),
    .A1(_20895_),
    .S(_00336_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _40921_ (.A0(_20895_),
    .A1(_00348_),
    .S(net101),
    .X(_00003_));
 sky130_fd_sc_hd__mux2_1 _40922_ (.A0(_02304_),
    .A1(_02305_),
    .S(\irq_state[1] ),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _40923_ (.A0(_02306_),
    .A1(_02304_),
    .S(_02217_),
    .X(_00008_));
 sky130_fd_sc_hd__mux2_1 _40924_ (.A0(_02214_),
    .A1(_02215_),
    .S(\irq_state[1] ),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _40925_ (.A0(_02216_),
    .A1(_02214_),
    .S(_02217_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _40926_ (.A0(_02218_),
    .A1(_02219_),
    .S(\irq_state[1] ),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _40927_ (.A0(_02220_),
    .A1(_02218_),
    .S(_02217_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _40928_ (.A0(_02221_),
    .A1(_02222_),
    .S(\irq_state[1] ),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _40929_ (.A0(_02223_),
    .A1(_02221_),
    .S(net424),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _40930_ (.A0(_02224_),
    .A1(_02225_),
    .S(\irq_state[1] ),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _40931_ (.A0(_02226_),
    .A1(_02224_),
    .S(net424),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _40932_ (.A0(_02227_),
    .A1(_02228_),
    .S(\irq_state[1] ),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _40933_ (.A0(_02229_),
    .A1(_02227_),
    .S(net424),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _40934_ (.A0(_02230_),
    .A1(_02231_),
    .S(\irq_state[1] ),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _40935_ (.A0(_02232_),
    .A1(_02230_),
    .S(net424),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _40936_ (.A0(_02233_),
    .A1(_02234_),
    .S(\irq_state[1] ),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _40937_ (.A0(_02235_),
    .A1(_02233_),
    .S(net424),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _40938_ (.A0(_02236_),
    .A1(_02237_),
    .S(\irq_state[1] ),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _40939_ (.A0(_02238_),
    .A1(_02236_),
    .S(net424),
    .X(_00009_));
 sky130_fd_sc_hd__mux2_1 _40940_ (.A0(_02239_),
    .A1(_02240_),
    .S(\irq_state[1] ),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _40941_ (.A0(_02241_),
    .A1(_02239_),
    .S(net424),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _40942_ (.A0(_02242_),
    .A1(_02243_),
    .S(\irq_state[1] ),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _40943_ (.A0(_02244_),
    .A1(_02242_),
    .S(net424),
    .X(_00011_));
 sky130_fd_sc_hd__mux2_1 _40944_ (.A0(_02245_),
    .A1(_02246_),
    .S(\irq_state[1] ),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _40945_ (.A0(_02247_),
    .A1(_02245_),
    .S(net424),
    .X(_00012_));
 sky130_fd_sc_hd__mux2_1 _40946_ (.A0(_02248_),
    .A1(_02249_),
    .S(\irq_state[1] ),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _40947_ (.A0(_02250_),
    .A1(_02248_),
    .S(net424),
    .X(_00013_));
 sky130_fd_sc_hd__mux2_1 _40948_ (.A0(_02251_),
    .A1(_02252_),
    .S(\irq_state[1] ),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _40949_ (.A0(_02253_),
    .A1(_02251_),
    .S(net424),
    .X(_00014_));
 sky130_fd_sc_hd__mux2_1 _40950_ (.A0(_02254_),
    .A1(_02255_),
    .S(\irq_state[1] ),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _40951_ (.A0(_02256_),
    .A1(_02254_),
    .S(net424),
    .X(_00015_));
 sky130_fd_sc_hd__mux2_1 _40952_ (.A0(_02257_),
    .A1(_02258_),
    .S(\irq_state[1] ),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _40953_ (.A0(_02259_),
    .A1(_02257_),
    .S(net424),
    .X(_00016_));
 sky130_fd_sc_hd__mux2_1 _40954_ (.A0(_02260_),
    .A1(_02261_),
    .S(\irq_state[1] ),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _40955_ (.A0(_02262_),
    .A1(_02260_),
    .S(net424),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _40956_ (.A0(_02263_),
    .A1(_02264_),
    .S(\irq_state[1] ),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _40957_ (.A0(_02265_),
    .A1(_02263_),
    .S(net424),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _40958_ (.A0(_02266_),
    .A1(_02267_),
    .S(\irq_state[1] ),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _40959_ (.A0(_02268_),
    .A1(_02266_),
    .S(net424),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _40960_ (.A0(_02269_),
    .A1(_02270_),
    .S(\irq_state[1] ),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _40961_ (.A0(_02271_),
    .A1(_02269_),
    .S(net424),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _40962_ (.A0(_02272_),
    .A1(_02273_),
    .S(\irq_state[1] ),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _40963_ (.A0(_02274_),
    .A1(_02272_),
    .S(net424),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _40964_ (.A0(_02275_),
    .A1(_02276_),
    .S(\irq_state[1] ),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _40965_ (.A0(_02277_),
    .A1(_02275_),
    .S(net424),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _40966_ (.A0(_02278_),
    .A1(_02279_),
    .S(\irq_state[1] ),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _40967_ (.A0(_02280_),
    .A1(_02278_),
    .S(net424),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _40968_ (.A0(_02281_),
    .A1(_02282_),
    .S(\irq_state[1] ),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _40969_ (.A0(_02283_),
    .A1(_02281_),
    .S(net424),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _40970_ (.A0(_02284_),
    .A1(_02285_),
    .S(\irq_state[1] ),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _40971_ (.A0(_02286_),
    .A1(_02284_),
    .S(net424),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _40972_ (.A0(_02287_),
    .A1(_02288_),
    .S(\irq_state[1] ),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _40973_ (.A0(_02289_),
    .A1(_02287_),
    .S(net424),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _40974_ (.A0(_02290_),
    .A1(_02291_),
    .S(\irq_state[1] ),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _40975_ (.A0(_02292_),
    .A1(_02290_),
    .S(net424),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _40976_ (.A0(_02293_),
    .A1(_02294_),
    .S(\irq_state[1] ),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _40977_ (.A0(_02295_),
    .A1(_02293_),
    .S(_02217_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _40978_ (.A0(_02296_),
    .A1(_02297_),
    .S(\irq_state[1] ),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _40979_ (.A0(_02298_),
    .A1(_02296_),
    .S(_02217_),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _40980_ (.A0(_02299_),
    .A1(_02300_),
    .S(\irq_state[1] ),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _40981_ (.A0(_02301_),
    .A1(_02299_),
    .S(_02217_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_2 _40982_ (.A0(_01467_),
    .A1(\reg_next_pc[1] ),
    .S(_00292_),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_2 _40983_ (.A0(_00295_),
    .A1(\reg_next_pc[2] ),
    .S(_00292_),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_2 _40984_ (.A0(_01470_),
    .A1(\reg_next_pc[3] ),
    .S(_00292_),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_2 _40985_ (.A0(_01478_),
    .A1(\reg_next_pc[5] ),
    .S(_00292_),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_2 _40986_ (.A0(_01481_),
    .A1(\reg_next_pc[6] ),
    .S(_00292_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_4 _40987_ (.A0(_01484_),
    .A1(\reg_next_pc[7] ),
    .S(_00292_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_2 _40988_ (.A0(_01487_),
    .A1(\reg_next_pc[8] ),
    .S(_00292_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_2 _40989_ (.A0(_01490_),
    .A1(\reg_next_pc[9] ),
    .S(_00292_),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_2 _40990_ (.A0(_01493_),
    .A1(\reg_next_pc[10] ),
    .S(_00292_),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_2 _40991_ (.A0(_01496_),
    .A1(\reg_next_pc[11] ),
    .S(_00292_),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_2 _40992_ (.A0(_01499_),
    .A1(\reg_next_pc[12] ),
    .S(_00292_),
    .X(_02561_));
 sky130_fd_sc_hd__mux2_2 _40993_ (.A0(_01502_),
    .A1(\reg_next_pc[13] ),
    .S(_00292_),
    .X(_02562_));
 sky130_fd_sc_hd__mux2_2 _40994_ (.A0(_01505_),
    .A1(\reg_next_pc[14] ),
    .S(_00292_),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_2 _40995_ (.A0(_01508_),
    .A1(\reg_next_pc[15] ),
    .S(_00292_),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_2 _40996_ (.A0(_01511_),
    .A1(\reg_next_pc[16] ),
    .S(_00292_),
    .X(_02565_));
 sky130_fd_sc_hd__mux2_2 _40997_ (.A0(_01514_),
    .A1(\reg_next_pc[17] ),
    .S(_00292_),
    .X(_02566_));
 sky130_fd_sc_hd__mux2_2 _40998_ (.A0(_01517_),
    .A1(\reg_next_pc[18] ),
    .S(_00292_),
    .X(_02567_));
 sky130_fd_sc_hd__mux2_2 _40999_ (.A0(_01520_),
    .A1(\reg_next_pc[19] ),
    .S(_00292_),
    .X(_02568_));
 sky130_fd_sc_hd__mux2_2 _41000_ (.A0(_01523_),
    .A1(\reg_next_pc[20] ),
    .S(_00292_),
    .X(_02569_));
 sky130_fd_sc_hd__mux2_4 _41001_ (.A0(_01526_),
    .A1(\reg_next_pc[21] ),
    .S(_00292_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_4 _41002_ (.A0(_01529_),
    .A1(\reg_next_pc[22] ),
    .S(_00292_),
    .X(_02572_));
 sky130_fd_sc_hd__mux2_2 _41003_ (.A0(_01532_),
    .A1(\reg_next_pc[23] ),
    .S(_00292_),
    .X(_02573_));
 sky130_fd_sc_hd__mux2_2 _41004_ (.A0(_01535_),
    .A1(\reg_next_pc[24] ),
    .S(_00292_),
    .X(_02574_));
 sky130_fd_sc_hd__mux2_4 _41005_ (.A0(_01538_),
    .A1(\reg_next_pc[25] ),
    .S(_00292_),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_4 _41006_ (.A0(_01541_),
    .A1(\reg_next_pc[26] ),
    .S(_00292_),
    .X(_02576_));
 sky130_fd_sc_hd__mux2_2 _41007_ (.A0(_01544_),
    .A1(\reg_next_pc[27] ),
    .S(_00292_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_2 _41008_ (.A0(_01547_),
    .A1(\reg_next_pc[28] ),
    .S(_00292_),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_2 _41009_ (.A0(_01550_),
    .A1(\reg_next_pc[29] ),
    .S(_00292_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_2 _41010_ (.A0(_01553_),
    .A1(\reg_next_pc[30] ),
    .S(_00292_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_2 _41011_ (.A0(_01556_),
    .A1(\reg_next_pc[31] ),
    .S(_00292_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _41012_ (.A0(_00057_),
    .A1(_00064_),
    .S(net225),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _41013_ (.A0(_00065_),
    .A1(_02543_),
    .S(net226),
    .X(_20931_));
 sky130_fd_sc_hd__mux2_1 _41014_ (.A0(_00075_),
    .A1(_00082_),
    .S(net503),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _41015_ (.A0(_00083_),
    .A1(_02544_),
    .S(net502),
    .X(_20932_));
 sky130_fd_sc_hd__mux2_1 _41016_ (.A0(_00089_),
    .A1(_00092_),
    .S(net503),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _41017_ (.A0(_00093_),
    .A1(_02545_),
    .S(net502),
    .X(_20933_));
 sky130_fd_sc_hd__mux2_1 _41018_ (.A0(_00099_),
    .A1(_00102_),
    .S(net503),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _41019_ (.A0(_00103_),
    .A1(_02546_),
    .S(net502),
    .X(_20934_));
 sky130_fd_sc_hd__mux2_1 _41020_ (.A0(_00107_),
    .A1(_00108_),
    .S(net225),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _41021_ (.A0(_00109_),
    .A1(_02547_),
    .S(net226),
    .X(_20935_));
 sky130_fd_sc_hd__mux2_1 _41022_ (.A0(_00113_),
    .A1(_00114_),
    .S(net503),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _41023_ (.A0(_00115_),
    .A1(_02548_),
    .S(net502),
    .X(_20936_));
 sky130_fd_sc_hd__mux2_1 _41024_ (.A0(_00119_),
    .A1(_00120_),
    .S(net225),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _41025_ (.A0(_00121_),
    .A1(_02549_),
    .S(net502),
    .X(_20937_));
 sky130_fd_sc_hd__mux2_1 _41026_ (.A0(_00125_),
    .A1(_00126_),
    .S(net503),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _41027_ (.A0(_00127_),
    .A1(_02550_),
    .S(net502),
    .X(_20938_));
 sky130_fd_sc_hd__mux2_1 _41028_ (.A0(_00129_),
    .A1(_00106_),
    .S(net222),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _41029_ (.A0(_00130_),
    .A1(_00057_),
    .S(net225),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _41030_ (.A0(_00131_),
    .A1(_02551_),
    .S(net226),
    .X(_20939_));
 sky130_fd_sc_hd__mux2_1 _41031_ (.A0(_00133_),
    .A1(_00112_),
    .S(net504),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _41032_ (.A0(_00134_),
    .A1(_00075_),
    .S(net503),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _41033_ (.A0(_00135_),
    .A1(_02552_),
    .S(net502),
    .X(_20940_));
 sky130_fd_sc_hd__mux2_1 _41034_ (.A0(_00137_),
    .A1(_00118_),
    .S(net222),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _41035_ (.A0(_00138_),
    .A1(_00089_),
    .S(net503),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _41036_ (.A0(_00139_),
    .A1(_02553_),
    .S(net502),
    .X(_20941_));
 sky130_fd_sc_hd__mux2_1 _41037_ (.A0(_00141_),
    .A1(_00124_),
    .S(net504),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _41038_ (.A0(_00142_),
    .A1(_00099_),
    .S(net503),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _41039_ (.A0(_00143_),
    .A1(_02554_),
    .S(net502),
    .X(_20942_));
 sky130_fd_sc_hd__mux2_1 _41040_ (.A0(_00144_),
    .A1(_00136_),
    .S(net211),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _41041_ (.A0(_00145_),
    .A1(_00129_),
    .S(net222),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _41042_ (.A0(_00146_),
    .A1(_00107_),
    .S(net225),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _41043_ (.A0(_00147_),
    .A1(_02555_),
    .S(net226),
    .X(_20943_));
 sky130_fd_sc_hd__mux2_1 _41044_ (.A0(_00148_),
    .A1(_00140_),
    .S(net505),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _41045_ (.A0(_00149_),
    .A1(_00133_),
    .S(net504),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _41046_ (.A0(_00150_),
    .A1(_00113_),
    .S(net503),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _41047_ (.A0(_00151_),
    .A1(_02556_),
    .S(net502),
    .X(_20944_));
 sky130_fd_sc_hd__mux2_1 _41048_ (.A0(net329),
    .A1(net327),
    .S(net200),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _41049_ (.A0(_00152_),
    .A1(_00144_),
    .S(net211),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _41050_ (.A0(_00153_),
    .A1(_00137_),
    .S(net222),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _41051_ (.A0(_00154_),
    .A1(_00119_),
    .S(net225),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _41052_ (.A0(_00155_),
    .A1(_02557_),
    .S(net226),
    .X(_20945_));
 sky130_fd_sc_hd__mux2_1 _41053_ (.A0(net330),
    .A1(net329),
    .S(net506),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _41054_ (.A0(_00156_),
    .A1(_00148_),
    .S(net505),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _41055_ (.A0(_00157_),
    .A1(_00141_),
    .S(net504),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _41056_ (.A0(_00158_),
    .A1(_00125_),
    .S(net503),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _41057_ (.A0(_00159_),
    .A1(_02558_),
    .S(net502),
    .X(_20946_));
 sky130_fd_sc_hd__mux2_1 _41058_ (.A0(net306),
    .A1(net317),
    .S(net506),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _41059_ (.A0(_00160_),
    .A1(_00161_),
    .S(net505),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _41060_ (.A0(_00162_),
    .A1(_00165_),
    .S(net504),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _41061_ (.A0(_00166_),
    .A1(_00173_),
    .S(net503),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _41062_ (.A0(_00174_),
    .A1(_00189_),
    .S(net502),
    .X(_20947_));
 sky130_fd_sc_hd__mux2_1 _41063_ (.A0(net317),
    .A1(net328),
    .S(net506),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _41064_ (.A0(_00190_),
    .A1(_00191_),
    .S(net505),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _41065_ (.A0(_00192_),
    .A1(_00195_),
    .S(net504),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _41066_ (.A0(_00196_),
    .A1(_00203_),
    .S(net503),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _41067_ (.A0(_00204_),
    .A1(_00220_),
    .S(net502),
    .X(_20958_));
 sky130_fd_sc_hd__mux2_1 _41068_ (.A0(_00161_),
    .A1(_00163_),
    .S(net505),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _41069_ (.A0(_00221_),
    .A1(_00222_),
    .S(net504),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _41070_ (.A0(_00223_),
    .A1(_00226_),
    .S(net503),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _41071_ (.A0(_00227_),
    .A1(_00234_),
    .S(net502),
    .X(_20969_));
 sky130_fd_sc_hd__mux2_1 _41072_ (.A0(_00191_),
    .A1(_00193_),
    .S(net505),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _41073_ (.A0(_00235_),
    .A1(_00236_),
    .S(net504),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _41074_ (.A0(_00237_),
    .A1(_00240_),
    .S(net503),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _41075_ (.A0(_00241_),
    .A1(_00248_),
    .S(net502),
    .X(_20972_));
 sky130_fd_sc_hd__mux2_1 _41076_ (.A0(_00165_),
    .A1(_00169_),
    .S(net504),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _41077_ (.A0(_00249_),
    .A1(_00250_),
    .S(net503),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _41078_ (.A0(_00251_),
    .A1(_00254_),
    .S(net502),
    .X(_20973_));
 sky130_fd_sc_hd__mux2_1 _41079_ (.A0(_00195_),
    .A1(_00199_),
    .S(net504),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _41080_ (.A0(_00255_),
    .A1(_00256_),
    .S(net503),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _41081_ (.A0(_00257_),
    .A1(_00260_),
    .S(net502),
    .X(_20974_));
 sky130_fd_sc_hd__mux2_1 _41082_ (.A0(_00222_),
    .A1(_00224_),
    .S(net504),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _41083_ (.A0(_00261_),
    .A1(_00262_),
    .S(net503),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _41084_ (.A0(_00263_),
    .A1(_00266_),
    .S(net502),
    .X(_20975_));
 sky130_fd_sc_hd__mux2_1 _41085_ (.A0(_00236_),
    .A1(_00238_),
    .S(net504),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _41086_ (.A0(_00267_),
    .A1(_00268_),
    .S(net503),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _41087_ (.A0(_00269_),
    .A1(_00272_),
    .S(net502),
    .X(_20976_));
 sky130_fd_sc_hd__mux2_1 _41088_ (.A0(_00173_),
    .A1(_00181_),
    .S(net503),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _41089_ (.A0(_00273_),
    .A1(_00274_),
    .S(net502),
    .X(_20977_));
 sky130_fd_sc_hd__mux2_1 _41090_ (.A0(_00203_),
    .A1(_00211_),
    .S(net503),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _41091_ (.A0(_00275_),
    .A1(_00276_),
    .S(net502),
    .X(_20978_));
 sky130_fd_sc_hd__mux2_1 _41092_ (.A0(_00226_),
    .A1(_00230_),
    .S(net503),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _41093_ (.A0(_00277_),
    .A1(_00278_),
    .S(net502),
    .X(_20948_));
 sky130_fd_sc_hd__mux2_1 _41094_ (.A0(_00240_),
    .A1(_00244_),
    .S(net503),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _41095_ (.A0(_00279_),
    .A1(_00280_),
    .S(net502),
    .X(_20949_));
 sky130_fd_sc_hd__mux2_1 _41096_ (.A0(_00250_),
    .A1(_00252_),
    .S(net503),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _41097_ (.A0(_00281_),
    .A1(_00282_),
    .S(net502),
    .X(_20950_));
 sky130_fd_sc_hd__mux2_1 _41098_ (.A0(_00256_),
    .A1(_00258_),
    .S(net503),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _41099_ (.A0(_00283_),
    .A1(_00284_),
    .S(net502),
    .X(_20951_));
 sky130_fd_sc_hd__mux2_1 _41100_ (.A0(_00262_),
    .A1(_00264_),
    .S(net503),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _41101_ (.A0(_00285_),
    .A1(_00286_),
    .S(net502),
    .X(_20952_));
 sky130_fd_sc_hd__mux2_1 _41102_ (.A0(_00268_),
    .A1(_00270_),
    .S(net503),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _41103_ (.A0(_00287_),
    .A1(_00288_),
    .S(net502),
    .X(_20953_));
 sky130_fd_sc_hd__mux2_1 _41104_ (.A0(_00189_),
    .A1(_00216_),
    .S(net502),
    .X(_20954_));
 sky130_fd_sc_hd__mux2_1 _41105_ (.A0(_00220_),
    .A1(_00216_),
    .S(net502),
    .X(_20955_));
 sky130_fd_sc_hd__mux2_1 _41106_ (.A0(_00234_),
    .A1(_00216_),
    .S(net502),
    .X(_20956_));
 sky130_fd_sc_hd__mux2_1 _41107_ (.A0(_00248_),
    .A1(_00216_),
    .S(net502),
    .X(_20957_));
 sky130_fd_sc_hd__mux2_1 _41108_ (.A0(_00254_),
    .A1(_00216_),
    .S(net502),
    .X(_20959_));
 sky130_fd_sc_hd__mux2_1 _41109_ (.A0(_00260_),
    .A1(_00216_),
    .S(net502),
    .X(_20960_));
 sky130_fd_sc_hd__mux2_1 _41110_ (.A0(_00266_),
    .A1(_00216_),
    .S(net502),
    .X(_20961_));
 sky130_fd_sc_hd__mux2_1 _41111_ (.A0(_00272_),
    .A1(_00216_),
    .S(net502),
    .X(_20962_));
 sky130_fd_sc_hd__mux2_1 _41112_ (.A0(_00274_),
    .A1(_00216_),
    .S(net502),
    .X(_20963_));
 sky130_fd_sc_hd__mux2_1 _41113_ (.A0(_00276_),
    .A1(_00216_),
    .S(net502),
    .X(_20964_));
 sky130_fd_sc_hd__mux2_1 _41114_ (.A0(_00278_),
    .A1(_00216_),
    .S(net502),
    .X(_20965_));
 sky130_fd_sc_hd__mux2_1 _41115_ (.A0(_00280_),
    .A1(_00216_),
    .S(net502),
    .X(_20966_));
 sky130_fd_sc_hd__mux2_1 _41116_ (.A0(_00282_),
    .A1(_00216_),
    .S(net502),
    .X(_20967_));
 sky130_fd_sc_hd__mux2_1 _41117_ (.A0(_00284_),
    .A1(_00216_),
    .S(net502),
    .X(_20968_));
 sky130_fd_sc_hd__mux2_1 _41118_ (.A0(_00286_),
    .A1(_00216_),
    .S(net502),
    .X(_20970_));
 sky130_fd_sc_hd__mux2_1 _41119_ (.A0(_00288_),
    .A1(_00216_),
    .S(net502),
    .X(_20971_));
 sky130_fd_sc_hd__mux2_1 _41120_ (.A0(_01697_),
    .A1(_01698_),
    .S(\irq_state[1] ),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _41121_ (.A0(_01705_),
    .A1(_01699_),
    .S(_01700_),
    .X(_20930_));
 sky130_fd_sc_hd__mux2_1 _41122_ (.A0(_01720_),
    .A1(\irq_pending[0] ),
    .S(_01706_),
    .X(_20896_));
 sky130_fd_sc_hd__mux2_1 _41123_ (.A0(_01733_),
    .A1(\irq_pending[1] ),
    .S(net464),
    .X(_20907_));
 sky130_fd_sc_hd__mux2_1 _41124_ (.A0(_01746_),
    .A1(\irq_pending[2] ),
    .S(net464),
    .X(_20918_));
 sky130_fd_sc_hd__mux2_1 _41125_ (.A0(_01759_),
    .A1(\irq_pending[3] ),
    .S(net464),
    .X(_20921_));
 sky130_fd_sc_hd__mux2_1 _41126_ (.A0(_01772_),
    .A1(\irq_pending[4] ),
    .S(net464),
    .X(_20922_));
 sky130_fd_sc_hd__mux2_1 _41127_ (.A0(_01785_),
    .A1(\irq_pending[5] ),
    .S(net464),
    .X(_20923_));
 sky130_fd_sc_hd__mux2_1 _41128_ (.A0(_01798_),
    .A1(\irq_pending[6] ),
    .S(net464),
    .X(_20924_));
 sky130_fd_sc_hd__mux2_1 _41129_ (.A0(_01811_),
    .A1(\irq_pending[7] ),
    .S(net464),
    .X(_20925_));
 sky130_fd_sc_hd__mux2_1 _41130_ (.A0(_01825_),
    .A1(\irq_pending[8] ),
    .S(net464),
    .X(_20926_));
 sky130_fd_sc_hd__mux2_1 _41131_ (.A0(_01838_),
    .A1(\irq_pending[9] ),
    .S(net463),
    .X(_20927_));
 sky130_fd_sc_hd__mux2_1 _41132_ (.A0(_01851_),
    .A1(\irq_pending[10] ),
    .S(net464),
    .X(_20897_));
 sky130_fd_sc_hd__mux2_1 _41133_ (.A0(_01864_),
    .A1(\irq_pending[11] ),
    .S(net464),
    .X(_20898_));
 sky130_fd_sc_hd__mux2_1 _41134_ (.A0(_01877_),
    .A1(\irq_pending[12] ),
    .S(net464),
    .X(_20899_));
 sky130_fd_sc_hd__mux2_1 _41135_ (.A0(_01890_),
    .A1(\irq_pending[13] ),
    .S(net464),
    .X(_20900_));
 sky130_fd_sc_hd__mux2_1 _41136_ (.A0(_01903_),
    .A1(\irq_pending[14] ),
    .S(net464),
    .X(_20901_));
 sky130_fd_sc_hd__mux2_1 _41137_ (.A0(_01916_),
    .A1(\irq_pending[15] ),
    .S(net464),
    .X(_20902_));
 sky130_fd_sc_hd__mux2_1 _41138_ (.A0(_01925_),
    .A1(\irq_pending[16] ),
    .S(net464),
    .X(_20903_));
 sky130_fd_sc_hd__mux2_1 _41139_ (.A0(_01934_),
    .A1(\irq_pending[17] ),
    .S(net463),
    .X(_20904_));
 sky130_fd_sc_hd__mux2_1 _41140_ (.A0(_01943_),
    .A1(\irq_pending[18] ),
    .S(net463),
    .X(_20905_));
 sky130_fd_sc_hd__mux2_1 _41141_ (.A0(_01952_),
    .A1(\irq_pending[19] ),
    .S(net463),
    .X(_20906_));
 sky130_fd_sc_hd__mux2_1 _41142_ (.A0(_01961_),
    .A1(\irq_pending[20] ),
    .S(net463),
    .X(_20908_));
 sky130_fd_sc_hd__mux2_1 _41143_ (.A0(_01970_),
    .A1(\irq_pending[21] ),
    .S(net463),
    .X(_20909_));
 sky130_fd_sc_hd__mux2_1 _41144_ (.A0(_01979_),
    .A1(\irq_pending[22] ),
    .S(net463),
    .X(_20910_));
 sky130_fd_sc_hd__mux2_1 _41145_ (.A0(_01988_),
    .A1(\irq_pending[23] ),
    .S(net463),
    .X(_20911_));
 sky130_fd_sc_hd__mux2_1 _41146_ (.A0(_01997_),
    .A1(\irq_pending[24] ),
    .S(net463),
    .X(_20912_));
 sky130_fd_sc_hd__mux2_1 _41147_ (.A0(_02006_),
    .A1(\irq_pending[25] ),
    .S(net463),
    .X(_20913_));
 sky130_fd_sc_hd__mux2_1 _41148_ (.A0(_02015_),
    .A1(\irq_pending[26] ),
    .S(net463),
    .X(_20914_));
 sky130_fd_sc_hd__mux2_1 _41149_ (.A0(_02024_),
    .A1(\irq_pending[27] ),
    .S(_01706_),
    .X(_20915_));
 sky130_fd_sc_hd__mux2_1 _41150_ (.A0(_02033_),
    .A1(\irq_pending[28] ),
    .S(_01706_),
    .X(_20916_));
 sky130_fd_sc_hd__mux2_1 _41151_ (.A0(_02042_),
    .A1(\irq_pending[29] ),
    .S(_01706_),
    .X(_20917_));
 sky130_fd_sc_hd__mux2_1 _41152_ (.A0(_02051_),
    .A1(\irq_pending[30] ),
    .S(_01706_),
    .X(_20919_));
 sky130_fd_sc_hd__mux2_1 _41153_ (.A0(_02060_),
    .A1(\irq_pending[31] ),
    .S(_01706_),
    .X(_20920_));
 sky130_fd_sc_hd__mux2_1 _41154_ (.A0(_02061_),
    .A1(net508),
    .S(_02542_),
    .X(_20891_));
 sky130_fd_sc_hd__mux2_4 _41155_ (.A0(\decoded_rd[0] ),
    .A1(\irq_state[0] ),
    .S(_00308_),
    .X(_20890_));
 sky130_fd_sc_hd__mux2_1 _41156_ (.A0(_02062_),
    .A1(_02065_),
    .S(_02542_),
    .X(_20928_));
 sky130_fd_sc_hd__mux2_1 _41157_ (.A0(_02068_),
    .A1(_02066_),
    .S(_02067_),
    .X(_20929_));
 sky130_fd_sc_hd__mux2_1 _41158_ (.A0(_02166_),
    .A1(_00291_),
    .S(_00290_),
    .X(_20892_));
 sky130_fd_sc_hd__mux2_1 _41159_ (.A0(_02166_),
    .A1(mem_do_wdata),
    .S(_00290_),
    .X(_20893_));
 sky130_fd_sc_hd__mux2_1 _41160_ (.A0(_00271_),
    .A1(_00216_),
    .S(net503),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _41161_ (.A0(_00265_),
    .A1(_00216_),
    .S(net503),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _41162_ (.A0(_00259_),
    .A1(_00216_),
    .S(net503),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _41163_ (.A0(_00253_),
    .A1(_00216_),
    .S(net503),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _41164_ (.A0(_00247_),
    .A1(_00216_),
    .S(net503),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _41165_ (.A0(_00233_),
    .A1(_00216_),
    .S(net503),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _41166_ (.A0(_00219_),
    .A1(_00216_),
    .S(net503),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _41167_ (.A0(_00188_),
    .A1(_00216_),
    .S(net503),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _41168_ (.A0(_00270_),
    .A1(_00271_),
    .S(net503),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _41169_ (.A0(_00246_),
    .A1(_00216_),
    .S(net504),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _41170_ (.A0(_00243_),
    .A1(_00245_),
    .S(net504),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _41171_ (.A0(_00239_),
    .A1(_00242_),
    .S(net504),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _41172_ (.A0(_00264_),
    .A1(_00265_),
    .S(net503),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _41173_ (.A0(_00232_),
    .A1(_00216_),
    .S(net504),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _41174_ (.A0(_00229_),
    .A1(_00231_),
    .S(net504),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _41175_ (.A0(_00225_),
    .A1(_00228_),
    .S(net504),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _41176_ (.A0(_00258_),
    .A1(_00259_),
    .S(net503),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _41177_ (.A0(_00218_),
    .A1(_00216_),
    .S(net504),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _41178_ (.A0(_00210_),
    .A1(_00214_),
    .S(net504),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _41179_ (.A0(_00202_),
    .A1(_00207_),
    .S(net504),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _41180_ (.A0(_00252_),
    .A1(_00253_),
    .S(net503),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _41181_ (.A0(_00187_),
    .A1(_00216_),
    .S(net504),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _41182_ (.A0(_00180_),
    .A1(_00184_),
    .S(net504),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _41183_ (.A0(_00172_),
    .A1(_00177_),
    .S(net504),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _41184_ (.A0(_00244_),
    .A1(_00247_),
    .S(net503),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _41185_ (.A0(_00245_),
    .A1(_00246_),
    .S(net504),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _41186_ (.A0(_00217_),
    .A1(_00216_),
    .S(net505),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _41187_ (.A0(_00213_),
    .A1(_00215_),
    .S(net505),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _41188_ (.A0(_00242_),
    .A1(_00243_),
    .S(net504),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _41189_ (.A0(_00209_),
    .A1(_00212_),
    .S(net505),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _41190_ (.A0(_00206_),
    .A1(_00208_),
    .S(net505),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _41191_ (.A0(_00238_),
    .A1(_00239_),
    .S(net504),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _41192_ (.A0(_00201_),
    .A1(_00205_),
    .S(net505),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _41193_ (.A0(_00198_),
    .A1(_00200_),
    .S(net505),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _41194_ (.A0(_00194_),
    .A1(_00197_),
    .S(net505),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _41195_ (.A0(_00230_),
    .A1(_00233_),
    .S(net503),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _41196_ (.A0(_00231_),
    .A1(_00232_),
    .S(net504),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _41197_ (.A0(_00186_),
    .A1(_00216_),
    .S(net505),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _41198_ (.A0(_00183_),
    .A1(_00185_),
    .S(net505),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _41199_ (.A0(_00228_),
    .A1(_00229_),
    .S(net504),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _41200_ (.A0(_00179_),
    .A1(_00182_),
    .S(net505),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _41201_ (.A0(_00176_),
    .A1(_00178_),
    .S(net505),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _41202_ (.A0(_00224_),
    .A1(_00225_),
    .S(net504),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _41203_ (.A0(_00171_),
    .A1(_00175_),
    .S(net505),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _41204_ (.A0(_00168_),
    .A1(_00170_),
    .S(net505),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _41205_ (.A0(_00164_),
    .A1(_00167_),
    .S(net505),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _41206_ (.A0(_00211_),
    .A1(_00219_),
    .S(net503),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _41207_ (.A0(_00214_),
    .A1(_00218_),
    .S(net504),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _41208_ (.A0(_00215_),
    .A1(_00217_),
    .S(net505),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _41209_ (.A0(net330),
    .A1(_00216_),
    .S(net506),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _41210_ (.A0(net327),
    .A1(net329),
    .S(net506),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _41211_ (.A0(_00212_),
    .A1(_00213_),
    .S(net505),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _41212_ (.A0(net325),
    .A1(net326),
    .S(net506),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _41213_ (.A0(net323),
    .A1(net324),
    .S(net506),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _41214_ (.A0(_00207_),
    .A1(_00210_),
    .S(net504),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _41215_ (.A0(_00208_),
    .A1(_00209_),
    .S(net505),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _41216_ (.A0(net321),
    .A1(net322),
    .S(net506),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _41217_ (.A0(net319),
    .A1(net320),
    .S(net506),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _41218_ (.A0(_00205_),
    .A1(_00206_),
    .S(net505),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _41219_ (.A0(net316),
    .A1(net318),
    .S(net506),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _41220_ (.A0(net314),
    .A1(net315),
    .S(net506),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _41221_ (.A0(_00199_),
    .A1(_00202_),
    .S(net504),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _41222_ (.A0(_00200_),
    .A1(_00201_),
    .S(net505),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _41223_ (.A0(net312),
    .A1(net313),
    .S(net506),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _41224_ (.A0(net310),
    .A1(net311),
    .S(net506),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _41225_ (.A0(_00197_),
    .A1(_00198_),
    .S(net505),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _41226_ (.A0(net308),
    .A1(net309),
    .S(net506),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _41227_ (.A0(net337),
    .A1(net307),
    .S(net506),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _41228_ (.A0(_00193_),
    .A1(_00194_),
    .S(net505),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _41229_ (.A0(net335),
    .A1(net336),
    .S(net506),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _41230_ (.A0(net333),
    .A1(net334),
    .S(net506),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _41231_ (.A0(net331),
    .A1(net332),
    .S(net506),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _41232_ (.A0(_00181_),
    .A1(_00188_),
    .S(net503),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _41233_ (.A0(_00184_),
    .A1(_00187_),
    .S(net504),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _41234_ (.A0(_00185_),
    .A1(_00186_),
    .S(net505),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _41235_ (.A0(net329),
    .A1(net330),
    .S(net506),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _41236_ (.A0(net326),
    .A1(net327),
    .S(net506),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _41237_ (.A0(_00182_),
    .A1(_00183_),
    .S(net505),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _41238_ (.A0(net324),
    .A1(net325),
    .S(net506),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _41239_ (.A0(net322),
    .A1(net323),
    .S(net506),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _41240_ (.A0(_00177_),
    .A1(_00180_),
    .S(net504),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _41241_ (.A0(_00178_),
    .A1(_00179_),
    .S(net505),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _41242_ (.A0(net320),
    .A1(net321),
    .S(net506),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _41243_ (.A0(net318),
    .A1(net319),
    .S(net506),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _41244_ (.A0(_00175_),
    .A1(_00176_),
    .S(net505),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _41245_ (.A0(net315),
    .A1(net316),
    .S(net506),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _41246_ (.A0(net313),
    .A1(net314),
    .S(net506),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _41247_ (.A0(_00169_),
    .A1(_00172_),
    .S(net504),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _41248_ (.A0(_00170_),
    .A1(_00171_),
    .S(net505),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _41249_ (.A0(net311),
    .A1(net312),
    .S(net506),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _41250_ (.A0(net309),
    .A1(net310),
    .S(net506),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _41251_ (.A0(_00167_),
    .A1(_00168_),
    .S(net505),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _41252_ (.A0(net307),
    .A1(net308),
    .S(net506),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _41253_ (.A0(net336),
    .A1(net337),
    .S(net506),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _41254_ (.A0(_00163_),
    .A1(_00164_),
    .S(net505),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _41255_ (.A0(net334),
    .A1(net335),
    .S(net506),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _41256_ (.A0(net332),
    .A1(net333),
    .S(net506),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _41257_ (.A0(net328),
    .A1(net331),
    .S(net506),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _41258_ (.A0(net327),
    .A1(net326),
    .S(net506),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _41259_ (.A0(net326),
    .A1(net325),
    .S(net200),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _41260_ (.A0(_00140_),
    .A1(_00132_),
    .S(net505),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _41261_ (.A0(net325),
    .A1(net324),
    .S(net506),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _41262_ (.A0(_00136_),
    .A1(_00128_),
    .S(net211),
    .X(_00137_));
 sky130_fd_sc_hd__mux2_1 _41263_ (.A0(net324),
    .A1(net323),
    .S(net200),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _41264_ (.A0(_00132_),
    .A1(_00123_),
    .S(net505),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _41265_ (.A0(net323),
    .A1(net322),
    .S(net506),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _41266_ (.A0(_00128_),
    .A1(_00117_),
    .S(net211),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _41267_ (.A0(net322),
    .A1(net321),
    .S(net200),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _41268_ (.A0(_00098_),
    .A1(_00100_),
    .S(net222),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _41269_ (.A0(_00124_),
    .A1(_00097_),
    .S(net504),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _41270_ (.A0(_00123_),
    .A1(_00111_),
    .S(net505),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _41271_ (.A0(net321),
    .A1(net320),
    .S(net506),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _41272_ (.A0(_00101_),
    .A1(_00094_),
    .S(net222),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _41273_ (.A0(_00088_),
    .A1(_00090_),
    .S(net222),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _41274_ (.A0(_00118_),
    .A1(_00087_),
    .S(net222),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _41275_ (.A0(_00117_),
    .A1(_00105_),
    .S(net211),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _41276_ (.A0(net320),
    .A1(net319),
    .S(net200),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _41277_ (.A0(_00091_),
    .A1(_00084_),
    .S(net222),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _41278_ (.A0(_00074_),
    .A1(_00078_),
    .S(net504),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _41279_ (.A0(_00112_),
    .A1(_00071_),
    .S(net504),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _41280_ (.A0(_00111_),
    .A1(_00096_),
    .S(net505),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _41281_ (.A0(net319),
    .A1(net318),
    .S(net506),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _41282_ (.A0(_00081_),
    .A1(_00067_),
    .S(net222),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _41283_ (.A0(_00056_),
    .A1(_00060_),
    .S(net222),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _41284_ (.A0(_00106_),
    .A1(_00053_),
    .S(net222),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _41285_ (.A0(_00105_),
    .A1(_00086_),
    .S(net211),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _41286_ (.A0(net318),
    .A1(net316),
    .S(net200),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _41287_ (.A0(_00063_),
    .A1(_00049_),
    .S(net222),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _41288_ (.A0(_00100_),
    .A1(_00101_),
    .S(net222),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _41289_ (.A0(_00077_),
    .A1(_00079_),
    .S(net505),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _41290_ (.A0(_00073_),
    .A1(_00076_),
    .S(net505),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _41291_ (.A0(_00097_),
    .A1(_00098_),
    .S(net504),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _41292_ (.A0(_00070_),
    .A1(_00072_),
    .S(net505),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _41293_ (.A0(_00096_),
    .A1(_00069_),
    .S(net505),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _41294_ (.A0(net316),
    .A1(net315),
    .S(net506),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _41295_ (.A0(_00080_),
    .A1(_00066_),
    .S(net505),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _41296_ (.A0(_00090_),
    .A1(_00091_),
    .S(net222),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _41297_ (.A0(_00059_),
    .A1(_00061_),
    .S(net211),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _41298_ (.A0(_00055_),
    .A1(_00058_),
    .S(net505),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _41299_ (.A0(_00087_),
    .A1(_00088_),
    .S(net222),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _41300_ (.A0(_00052_),
    .A1(_00054_),
    .S(net211),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _41301_ (.A0(_00086_),
    .A1(_00051_),
    .S(net211),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _41302_ (.A0(net315),
    .A1(net314),
    .S(net200),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_2 _41303_ (.A0(_00062_),
    .A1(_00048_),
    .S(net211),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _41304_ (.A0(_00078_),
    .A1(_00081_),
    .S(net504),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _41305_ (.A0(_00079_),
    .A1(_00080_),
    .S(net505),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _41306_ (.A0(net331),
    .A1(net328),
    .S(net200),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _41307_ (.A0(net333),
    .A1(net332),
    .S(net200),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _41308_ (.A0(_00076_),
    .A1(_00077_),
    .S(net505),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _41309_ (.A0(net335),
    .A1(net334),
    .S(net200),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _41310_ (.A0(net337),
    .A1(net336),
    .S(net200),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _41311_ (.A0(_00071_),
    .A1(_00074_),
    .S(net504),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _41312_ (.A0(_00072_),
    .A1(_00073_),
    .S(net505),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _41313_ (.A0(net308),
    .A1(net307),
    .S(net506),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _41314_ (.A0(net310),
    .A1(net309),
    .S(net506),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _41315_ (.A0(_00069_),
    .A1(_00070_),
    .S(net505),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _41316_ (.A0(net312),
    .A1(net311),
    .S(net506),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _41317_ (.A0(net314),
    .A1(net313),
    .S(net506),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _41318_ (.A0(net317),
    .A1(net306),
    .S(net200),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _41319_ (.A0(_00060_),
    .A1(_00063_),
    .S(net222),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _41320_ (.A0(_00061_),
    .A1(_00062_),
    .S(net211),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _41321_ (.A0(net328),
    .A1(net317),
    .S(net200),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _41322_ (.A0(net332),
    .A1(net331),
    .S(net200),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _41323_ (.A0(_00058_),
    .A1(_00059_),
    .S(net211),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _41324_ (.A0(net334),
    .A1(net333),
    .S(net200),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _41325_ (.A0(net336),
    .A1(net335),
    .S(net200),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _41326_ (.A0(_00053_),
    .A1(_00056_),
    .S(net222),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _41327_ (.A0(_00054_),
    .A1(_00055_),
    .S(net211),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _41328_ (.A0(net307),
    .A1(net337),
    .S(net200),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _41329_ (.A0(net309),
    .A1(net308),
    .S(net506),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _41330_ (.A0(_00051_),
    .A1(_00052_),
    .S(net211),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _41331_ (.A0(net311),
    .A1(net310),
    .S(net200),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _41332_ (.A0(net313),
    .A1(net312),
    .S(net506),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _41333_ (.A0(_02408_),
    .A1(net362),
    .S(instr_sub),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_2 _41334_ (.A0(_02406_),
    .A1(_02405_),
    .S(instr_sub),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_2 _41335_ (.A0(_02403_),
    .A1(_02402_),
    .S(instr_sub),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _41336_ (.A0(_02400_),
    .A1(_02399_),
    .S(instr_sub),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _41337_ (.A0(_02397_),
    .A1(_02396_),
    .S(instr_sub),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _41338_ (.A0(_02394_),
    .A1(_02393_),
    .S(instr_sub),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _41339_ (.A0(_02391_),
    .A1(_02390_),
    .S(instr_sub),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _41340_ (.A0(_02388_),
    .A1(_02387_),
    .S(instr_sub),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _41341_ (.A0(_02385_),
    .A1(_02384_),
    .S(instr_sub),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _41342_ (.A0(_02382_),
    .A1(_02381_),
    .S(instr_sub),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_2 _41343_ (.A0(_02379_),
    .A1(_02378_),
    .S(instr_sub),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_2 _41344_ (.A0(_02376_),
    .A1(_02375_),
    .S(instr_sub),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_2 _41345_ (.A0(_02373_),
    .A1(_02372_),
    .S(instr_sub),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_2 _41346_ (.A0(_02370_),
    .A1(_02369_),
    .S(instr_sub),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _41347_ (.A0(_02367_),
    .A1(_02366_),
    .S(instr_sub),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_2 _41348_ (.A0(_02364_),
    .A1(_02363_),
    .S(instr_sub),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _41349_ (.A0(_02361_),
    .A1(_02360_),
    .S(instr_sub),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _41350_ (.A0(_02358_),
    .A1(_02357_),
    .S(instr_sub),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _41351_ (.A0(_02355_),
    .A1(_02354_),
    .S(instr_sub),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _41352_ (.A0(_02352_),
    .A1(_02351_),
    .S(instr_sub),
    .X(_02353_));
 sky130_fd_sc_hd__mux2_1 _41353_ (.A0(_02349_),
    .A1(_02348_),
    .S(instr_sub),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _41354_ (.A0(_02346_),
    .A1(_02345_),
    .S(instr_sub),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _41355_ (.A0(_02343_),
    .A1(_02342_),
    .S(instr_sub),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _41356_ (.A0(_02340_),
    .A1(_02339_),
    .S(instr_sub),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _41357_ (.A0(_02337_),
    .A1(_02336_),
    .S(instr_sub),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_4 _41358_ (.A0(_02334_),
    .A1(_02333_),
    .S(instr_sub),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _41359_ (.A0(_02331_),
    .A1(_02330_),
    .S(instr_sub),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _41360_ (.A0(_02328_),
    .A1(_02327_),
    .S(instr_sub),
    .X(_02329_));
 sky130_fd_sc_hd__mux2_1 _41361_ (.A0(_02325_),
    .A1(_02324_),
    .S(instr_sub),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _41362_ (.A0(_02322_),
    .A1(_02321_),
    .S(instr_sub),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _41363_ (.A0(_02319_),
    .A1(_02318_),
    .S(instr_sub),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _41364_ (.A0(_02313_),
    .A1(_02314_),
    .S(_00306_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _41365_ (.A0(_02311_),
    .A1(_02315_),
    .S(_00303_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _41366_ (.A0(_02311_),
    .A1(_02312_),
    .S(_00305_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _41367_ (.A0(_02307_),
    .A1(_02308_),
    .S(\irq_state[1] ),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _41368_ (.A0(_02309_),
    .A1(_02307_),
    .S(_02217_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _41369_ (.A0(_02302_),
    .A1(\irq_pending[0] ),
    .S(_01208_),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _41370_ (.A0(\reg_out[0] ),
    .A1(\alu_out_q[0] ),
    .S(latched_stalu),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _41371_ (.A0(_02063_),
    .A1(_00343_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _41372_ (.A0(_02056_),
    .A1(_02055_),
    .S(_01714_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_2 _41373_ (.A0(_02058_),
    .A1(_02057_),
    .S(_01717_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_2 _41374_ (.A0(\pcpi_mul.rd[31] ),
    .A1(\pcpi_mul.rd[63] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _41375_ (.A0(_01908_),
    .A1(_02052_),
    .S(net496),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _41376_ (.A0(_02047_),
    .A1(_02046_),
    .S(_01714_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_2 _41377_ (.A0(_02049_),
    .A1(_02048_),
    .S(_01717_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_2 _41378_ (.A0(\pcpi_mul.rd[30] ),
    .A1(\pcpi_mul.rd[62] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _41379_ (.A0(_01908_),
    .A1(_02043_),
    .S(net496),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _41380_ (.A0(_02038_),
    .A1(_02037_),
    .S(_01714_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_2 _41381_ (.A0(_02040_),
    .A1(_02039_),
    .S(_01717_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _41382_ (.A0(\pcpi_mul.rd[29] ),
    .A1(\pcpi_mul.rd[61] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _41383_ (.A0(_01908_),
    .A1(_02034_),
    .S(net496),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _41384_ (.A0(_02029_),
    .A1(_02028_),
    .S(_01714_),
    .X(_02030_));
 sky130_fd_sc_hd__mux2_2 _41385_ (.A0(_02031_),
    .A1(_02030_),
    .S(_01717_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_2 _41386_ (.A0(\pcpi_mul.rd[28] ),
    .A1(\pcpi_mul.rd[60] ),
    .S(\pcpi_mul.shift_out ),
    .X(_02027_));
 sky130_fd_sc_hd__mux2_1 _41387_ (.A0(_01908_),
    .A1(_02025_),
    .S(net496),
    .X(_02026_));
 sky130_fd_sc_hd__mux2_1 _41388_ (.A0(_02020_),
    .A1(_02019_),
    .S(_01714_),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_2 _41389_ (.A0(_02022_),
    .A1(_02021_),
    .S(_01717_),
    .X(_02023_));
 sky130_fd_sc_hd__mux2_1 _41390_ (.A0(\pcpi_mul.rd[27] ),
    .A1(\pcpi_mul.rd[59] ),
    .S(net509),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _41391_ (.A0(_01908_),
    .A1(_02016_),
    .S(net496),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _41392_ (.A0(_02011_),
    .A1(_02010_),
    .S(_01714_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_2 _41393_ (.A0(_02013_),
    .A1(_02012_),
    .S(_01717_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _41394_ (.A0(\pcpi_mul.rd[26] ),
    .A1(\pcpi_mul.rd[58] ),
    .S(net509),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _41395_ (.A0(_01908_),
    .A1(_02007_),
    .S(net496),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _41396_ (.A0(_02002_),
    .A1(_02001_),
    .S(_01714_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_2 _41397_ (.A0(_02004_),
    .A1(_02003_),
    .S(_01717_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _41398_ (.A0(\pcpi_mul.rd[25] ),
    .A1(\pcpi_mul.rd[57] ),
    .S(net509),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _41399_ (.A0(_01908_),
    .A1(_01998_),
    .S(net496),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _41400_ (.A0(_01993_),
    .A1(_01992_),
    .S(_01714_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _41401_ (.A0(_01995_),
    .A1(_01994_),
    .S(_01717_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _41402_ (.A0(\pcpi_mul.rd[24] ),
    .A1(\pcpi_mul.rd[56] ),
    .S(net509),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_2 _41403_ (.A0(_01908_),
    .A1(_01989_),
    .S(net496),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_2 _41404_ (.A0(_01984_),
    .A1(_01983_),
    .S(_01714_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_2 _41405_ (.A0(_01986_),
    .A1(_01985_),
    .S(_01717_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _41406_ (.A0(\pcpi_mul.rd[23] ),
    .A1(\pcpi_mul.rd[55] ),
    .S(net509),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _41407_ (.A0(_01908_),
    .A1(_01980_),
    .S(net496),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _41408_ (.A0(_01975_),
    .A1(_01974_),
    .S(_01714_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_2 _41409_ (.A0(_01977_),
    .A1(_01976_),
    .S(_01717_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _41410_ (.A0(\pcpi_mul.rd[22] ),
    .A1(\pcpi_mul.rd[54] ),
    .S(net509),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _41411_ (.A0(_01908_),
    .A1(_01971_),
    .S(net496),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_2 _41412_ (.A0(_01966_),
    .A1(_01965_),
    .S(_01714_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_2 _41413_ (.A0(_01968_),
    .A1(_01967_),
    .S(_01717_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _41414_ (.A0(\pcpi_mul.rd[21] ),
    .A1(\pcpi_mul.rd[53] ),
    .S(net509),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _41415_ (.A0(_01908_),
    .A1(_01962_),
    .S(net496),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_2 _41416_ (.A0(_01957_),
    .A1(_01956_),
    .S(_01714_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_2 _41417_ (.A0(_01959_),
    .A1(_01958_),
    .S(_01717_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _41418_ (.A0(\pcpi_mul.rd[20] ),
    .A1(\pcpi_mul.rd[52] ),
    .S(\pcpi_mul.shift_out ),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _41419_ (.A0(_01908_),
    .A1(_01953_),
    .S(net496),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_2 _41420_ (.A0(_01948_),
    .A1(_01947_),
    .S(_01714_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_2 _41421_ (.A0(_01950_),
    .A1(_01949_),
    .S(_01717_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _41422_ (.A0(\pcpi_mul.rd[19] ),
    .A1(\pcpi_mul.rd[51] ),
    .S(net509),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _41423_ (.A0(_01908_),
    .A1(_01944_),
    .S(net496),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _41424_ (.A0(_01939_),
    .A1(_01938_),
    .S(_01714_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_2 _41425_ (.A0(_01941_),
    .A1(_01940_),
    .S(_01717_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _41426_ (.A0(\pcpi_mul.rd[18] ),
    .A1(\pcpi_mul.rd[50] ),
    .S(net509),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _41427_ (.A0(_01908_),
    .A1(_01935_),
    .S(net496),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_2 _41428_ (.A0(_01930_),
    .A1(_01929_),
    .S(_01714_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_2 _41429_ (.A0(_01932_),
    .A1(_01931_),
    .S(_01717_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _41430_ (.A0(\pcpi_mul.rd[17] ),
    .A1(\pcpi_mul.rd[49] ),
    .S(net509),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _41431_ (.A0(_01908_),
    .A1(_01926_),
    .S(net496),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _41432_ (.A0(_01921_),
    .A1(_01920_),
    .S(_01714_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_2 _41433_ (.A0(_01923_),
    .A1(_01922_),
    .S(_01717_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _41434_ (.A0(\pcpi_mul.rd[16] ),
    .A1(\pcpi_mul.rd[48] ),
    .S(net509),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _41435_ (.A0(_01908_),
    .A1(_01917_),
    .S(net496),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_2 _41436_ (.A0(_01912_),
    .A1(_01911_),
    .S(_01714_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_2 _41437_ (.A0(_01914_),
    .A1(_01913_),
    .S(_01717_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _41438_ (.A0(\pcpi_mul.rd[15] ),
    .A1(\pcpi_mul.rd[47] ),
    .S(net509),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_2 _41439_ (.A0(_01908_),
    .A1(_01907_),
    .S(net496),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_2 _41440_ (.A0(_01906_),
    .A1(_01904_),
    .S(net431),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _41441_ (.A0(net516),
    .A1(net57),
    .S(net317),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_2 _41442_ (.A0(_01899_),
    .A1(_01898_),
    .S(_01714_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_2 _41443_ (.A0(_01901_),
    .A1(_01900_),
    .S(_01717_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _41444_ (.A0(\pcpi_mul.rd[14] ),
    .A1(\pcpi_mul.rd[46] ),
    .S(net509),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_2 _41445_ (.A0(_01895_),
    .A1(_01894_),
    .S(net496),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _41446_ (.A0(_01893_),
    .A1(_01891_),
    .S(net431),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _41447_ (.A0(net38),
    .A1(net513),
    .S(net317),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _41448_ (.A0(_01886_),
    .A1(_01885_),
    .S(_01714_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_2 _41449_ (.A0(_01888_),
    .A1(_01887_),
    .S(_01717_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _41450_ (.A0(\pcpi_mul.rd[13] ),
    .A1(\pcpi_mul.rd[45] ),
    .S(net509),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _41451_ (.A0(_01882_),
    .A1(_01881_),
    .S(_01816_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _41452_ (.A0(_01880_),
    .A1(_01878_),
    .S(net431),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _41453_ (.A0(net37),
    .A1(net54),
    .S(net317),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_2 _41454_ (.A0(_01873_),
    .A1(_01872_),
    .S(_01714_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_2 _41455_ (.A0(_01875_),
    .A1(_01874_),
    .S(_01717_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _41456_ (.A0(\pcpi_mul.rd[12] ),
    .A1(\pcpi_mul.rd[44] ),
    .S(net509),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_2 _41457_ (.A0(_01869_),
    .A1(_01868_),
    .S(_01816_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _41458_ (.A0(_01867_),
    .A1(_01865_),
    .S(net431),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _41459_ (.A0(net517),
    .A1(net53),
    .S(net317),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_2 _41460_ (.A0(_01860_),
    .A1(_01859_),
    .S(_01714_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_2 _41461_ (.A0(_01862_),
    .A1(_01861_),
    .S(_01717_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_4 _41462_ (.A0(\pcpi_mul.rd[11] ),
    .A1(\pcpi_mul.rd[43] ),
    .S(net509),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _41463_ (.A0(_01856_),
    .A1(_01855_),
    .S(_01816_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _41464_ (.A0(_01854_),
    .A1(_01852_),
    .S(net431),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _41465_ (.A0(net35),
    .A1(net52),
    .S(net317),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_2 _41466_ (.A0(_01847_),
    .A1(_01846_),
    .S(_01714_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_2 _41467_ (.A0(_01849_),
    .A1(_01848_),
    .S(_01717_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_4 _41468_ (.A0(\pcpi_mul.rd[10] ),
    .A1(\pcpi_mul.rd[42] ),
    .S(net509),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_2 _41469_ (.A0(_01843_),
    .A1(_01842_),
    .S(_01816_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _41470_ (.A0(_01841_),
    .A1(_01839_),
    .S(net431),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _41471_ (.A0(net34),
    .A1(net51),
    .S(net317),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_4 _41472_ (.A0(_01834_),
    .A1(_01833_),
    .S(_01714_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _41473_ (.A0(_01836_),
    .A1(_01835_),
    .S(_01717_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_4 _41474_ (.A0(\pcpi_mul.rd[9] ),
    .A1(\pcpi_mul.rd[41] ),
    .S(net509),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_2 _41475_ (.A0(_01830_),
    .A1(_01829_),
    .S(_01816_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _41476_ (.A0(_01828_),
    .A1(_01826_),
    .S(net431),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _41477_ (.A0(net64),
    .A1(net50),
    .S(net317),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_4 _41478_ (.A0(_01821_),
    .A1(_01820_),
    .S(_01714_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_2 _41479_ (.A0(_01823_),
    .A1(_01822_),
    .S(_01717_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_4 _41480_ (.A0(\pcpi_mul.rd[8] ),
    .A1(\pcpi_mul.rd[40] ),
    .S(net509),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_2 _41481_ (.A0(_01817_),
    .A1(_01815_),
    .S(_01816_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _41482_ (.A0(_01814_),
    .A1(_01812_),
    .S(net431),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _41483_ (.A0(net63),
    .A1(net49),
    .S(net317),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_2 _41484_ (.A0(_01807_),
    .A1(_01806_),
    .S(_01714_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _41485_ (.A0(_01809_),
    .A1(_01808_),
    .S(_01717_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_4 _41486_ (.A0(\pcpi_mul.rd[7] ),
    .A1(\pcpi_mul.rd[39] ),
    .S(net509),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _41487_ (.A0(_01803_),
    .A1(_01799_),
    .S(net431),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _41488_ (.A0(net62),
    .A1(net48),
    .S(net317),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _41489_ (.A0(_01800_),
    .A1(_01799_),
    .S(_00304_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_2 _41490_ (.A0(_01794_),
    .A1(_01793_),
    .S(_01714_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_2 _41491_ (.A0(_01796_),
    .A1(_01795_),
    .S(_01717_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_4 _41492_ (.A0(\pcpi_mul.rd[6] ),
    .A1(\pcpi_mul.rd[38] ),
    .S(net509),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_2 _41493_ (.A0(_01790_),
    .A1(_01786_),
    .S(net431),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _41494_ (.A0(net61),
    .A1(net47),
    .S(net317),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _41495_ (.A0(_01787_),
    .A1(_01786_),
    .S(_00304_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_2 _41496_ (.A0(_01781_),
    .A1(_01780_),
    .S(_01714_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _41497_ (.A0(_01783_),
    .A1(_01782_),
    .S(_01717_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_4 _41498_ (.A0(\pcpi_mul.rd[5] ),
    .A1(\pcpi_mul.rd[37] ),
    .S(net509),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_2 _41499_ (.A0(_01777_),
    .A1(_01773_),
    .S(net431),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _41500_ (.A0(net512),
    .A1(net46),
    .S(net317),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _41501_ (.A0(_01774_),
    .A1(_01773_),
    .S(_00304_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_2 _41502_ (.A0(_01768_),
    .A1(_01767_),
    .S(_01714_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_2 _41503_ (.A0(_01770_),
    .A1(_01769_),
    .S(_01717_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_4 _41504_ (.A0(\pcpi_mul.rd[4] ),
    .A1(\pcpi_mul.rd[36] ),
    .S(net509),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_2 _41505_ (.A0(_01764_),
    .A1(_01760_),
    .S(net431),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _41506_ (.A0(net59),
    .A1(net514),
    .S(net317),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _41507_ (.A0(_01761_),
    .A1(_01760_),
    .S(_00304_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_2 _41508_ (.A0(_01755_),
    .A1(_01754_),
    .S(_01714_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _41509_ (.A0(_01757_),
    .A1(_01756_),
    .S(_01717_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_4 _41510_ (.A0(\pcpi_mul.rd[3] ),
    .A1(\pcpi_mul.rd[35] ),
    .S(net509),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _41511_ (.A0(_01751_),
    .A1(_01747_),
    .S(net431),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _41512_ (.A0(net58),
    .A1(net515),
    .S(net317),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _41513_ (.A0(_01748_),
    .A1(_01747_),
    .S(_00304_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_2 _41514_ (.A0(_01742_),
    .A1(_01741_),
    .S(_01714_),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _41515_ (.A0(_01744_),
    .A1(_01743_),
    .S(_01717_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_4 _41516_ (.A0(\pcpi_mul.rd[2] ),
    .A1(\pcpi_mul.rd[34] ),
    .S(net509),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _41517_ (.A0(_01738_),
    .A1(_01734_),
    .S(net431),
    .X(_01739_));
 sky130_fd_sc_hd__mux2_1 _41518_ (.A0(net55),
    .A1(net42),
    .S(net317),
    .X(_01737_));
 sky130_fd_sc_hd__mux2_1 _41519_ (.A0(_01735_),
    .A1(_01734_),
    .S(_00304_),
    .X(_01736_));
 sky130_fd_sc_hd__mux2_2 _41520_ (.A0(_01729_),
    .A1(_01728_),
    .S(_01714_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _41521_ (.A0(_01731_),
    .A1(_01730_),
    .S(_01717_),
    .X(_01732_));
 sky130_fd_sc_hd__mux2_1 _41522_ (.A0(\pcpi_mul.rd[1] ),
    .A1(\pcpi_mul.rd[33] ),
    .S(net509),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _41523_ (.A0(_01725_),
    .A1(_01721_),
    .S(net431),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _41524_ (.A0(net44),
    .A1(net41),
    .S(net317),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _41525_ (.A0(_01722_),
    .A1(_01721_),
    .S(_00304_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_2 _41526_ (.A0(_01715_),
    .A1(_02559_),
    .S(_01714_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_2 _41527_ (.A0(_01718_),
    .A1(_01716_),
    .S(_01717_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_2 _41528_ (.A0(\pcpi_mul.rd[0] ),
    .A1(\pcpi_mul.rd[32] ),
    .S(net509),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _41529_ (.A0(_01711_),
    .A1(_01707_),
    .S(net431),
    .X(_01712_));
 sky130_fd_sc_hd__mux2_1 _41530_ (.A0(net33),
    .A1(net40),
    .S(net317),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _41531_ (.A0(_01708_),
    .A1(_01707_),
    .S(_00304_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _41532_ (.A0(_01701_),
    .A1(_01696_),
    .S(_00311_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _41533_ (.A0(_01702_),
    .A1(_01696_),
    .S(\pcpi_mul.active[1] ),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _41534_ (.A0(_01696_),
    .A1(_01703_),
    .S(_00310_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _41535_ (.A0(_01693_),
    .A1(net273),
    .S(_00316_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _41536_ (.A0(_01690_),
    .A1(net272),
    .S(_00316_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _41537_ (.A0(_01687_),
    .A1(net271),
    .S(_00316_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _41538_ (.A0(_01684_),
    .A1(net270),
    .S(_00316_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _41539_ (.A0(\reg_next_pc[31] ),
    .A1(_01554_),
    .S(latched_store),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _41540_ (.A0(\reg_out[31] ),
    .A1(\alu_out_q[31] ),
    .S(latched_stalu),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _41541_ (.A0(\reg_next_pc[30] ),
    .A1(_01551_),
    .S(latched_store),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_2 _41542_ (.A0(\reg_out[30] ),
    .A1(\alu_out_q[30] ),
    .S(latched_stalu),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _41543_ (.A0(\reg_next_pc[29] ),
    .A1(_01548_),
    .S(latched_store),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_2 _41544_ (.A0(\reg_out[29] ),
    .A1(\alu_out_q[29] ),
    .S(latched_stalu),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _41545_ (.A0(\reg_next_pc[28] ),
    .A1(_01545_),
    .S(latched_store),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_2 _41546_ (.A0(\reg_out[28] ),
    .A1(\alu_out_q[28] ),
    .S(latched_stalu),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _41547_ (.A0(\reg_next_pc[27] ),
    .A1(_01542_),
    .S(latched_store),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_2 _41548_ (.A0(\reg_out[27] ),
    .A1(\alu_out_q[27] ),
    .S(latched_stalu),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _41549_ (.A0(\reg_next_pc[26] ),
    .A1(_01539_),
    .S(latched_store),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _41550_ (.A0(\reg_out[26] ),
    .A1(\alu_out_q[26] ),
    .S(latched_stalu),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _41551_ (.A0(\reg_next_pc[25] ),
    .A1(_01536_),
    .S(latched_store),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _41552_ (.A0(\reg_out[25] ),
    .A1(\alu_out_q[25] ),
    .S(latched_stalu),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _41553_ (.A0(\reg_next_pc[24] ),
    .A1(_01533_),
    .S(latched_store),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _41554_ (.A0(\reg_out[24] ),
    .A1(\alu_out_q[24] ),
    .S(latched_stalu),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _41555_ (.A0(\reg_next_pc[23] ),
    .A1(_01530_),
    .S(latched_store),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _41556_ (.A0(\reg_out[23] ),
    .A1(\alu_out_q[23] ),
    .S(latched_stalu),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _41557_ (.A0(\reg_next_pc[22] ),
    .A1(_01527_),
    .S(latched_store),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _41558_ (.A0(\reg_out[22] ),
    .A1(\alu_out_q[22] ),
    .S(latched_stalu),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _41559_ (.A0(\reg_next_pc[21] ),
    .A1(_01524_),
    .S(latched_store),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _41560_ (.A0(\reg_out[21] ),
    .A1(\alu_out_q[21] ),
    .S(latched_stalu),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _41561_ (.A0(\reg_next_pc[20] ),
    .A1(_01521_),
    .S(latched_store),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _41562_ (.A0(\reg_out[20] ),
    .A1(\alu_out_q[20] ),
    .S(latched_stalu),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _41563_ (.A0(\reg_next_pc[19] ),
    .A1(_01518_),
    .S(latched_store),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _41564_ (.A0(\reg_out[19] ),
    .A1(\alu_out_q[19] ),
    .S(latched_stalu),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _41565_ (.A0(\reg_next_pc[18] ),
    .A1(_01515_),
    .S(latched_store),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _41566_ (.A0(\reg_out[18] ),
    .A1(\alu_out_q[18] ),
    .S(latched_stalu),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _41567_ (.A0(\reg_next_pc[17] ),
    .A1(_01512_),
    .S(latched_store),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _41568_ (.A0(\reg_out[17] ),
    .A1(\alu_out_q[17] ),
    .S(latched_stalu),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _41569_ (.A0(\reg_next_pc[16] ),
    .A1(_01509_),
    .S(latched_store),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _41570_ (.A0(\reg_out[16] ),
    .A1(\alu_out_q[16] ),
    .S(latched_stalu),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _41571_ (.A0(\reg_next_pc[15] ),
    .A1(_01506_),
    .S(latched_store),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _41572_ (.A0(\reg_out[15] ),
    .A1(\alu_out_q[15] ),
    .S(latched_stalu),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _41573_ (.A0(\reg_next_pc[14] ),
    .A1(_01503_),
    .S(latched_store),
    .X(_01504_));
 sky130_fd_sc_hd__mux2_1 _41574_ (.A0(\reg_out[14] ),
    .A1(\alu_out_q[14] ),
    .S(latched_stalu),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _41575_ (.A0(\reg_next_pc[13] ),
    .A1(_01500_),
    .S(latched_store),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_2 _41576_ (.A0(\reg_out[13] ),
    .A1(\alu_out_q[13] ),
    .S(latched_stalu),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _41577_ (.A0(\reg_next_pc[12] ),
    .A1(_01497_),
    .S(latched_store),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _41578_ (.A0(\reg_out[12] ),
    .A1(\alu_out_q[12] ),
    .S(latched_stalu),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _41579_ (.A0(\reg_next_pc[11] ),
    .A1(_01494_),
    .S(latched_store),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _41580_ (.A0(\reg_out[11] ),
    .A1(\alu_out_q[11] ),
    .S(latched_stalu),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _41581_ (.A0(\reg_next_pc[10] ),
    .A1(_01491_),
    .S(latched_store),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _41582_ (.A0(\reg_out[10] ),
    .A1(\alu_out_q[10] ),
    .S(latched_stalu),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _41583_ (.A0(\reg_next_pc[9] ),
    .A1(_01488_),
    .S(latched_store),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _41584_ (.A0(\reg_out[9] ),
    .A1(\alu_out_q[9] ),
    .S(latched_stalu),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _41585_ (.A0(\reg_next_pc[8] ),
    .A1(_01485_),
    .S(latched_store),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _41586_ (.A0(\reg_out[8] ),
    .A1(\alu_out_q[8] ),
    .S(latched_stalu),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _41587_ (.A0(\reg_next_pc[7] ),
    .A1(_01482_),
    .S(latched_store),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _41588_ (.A0(\reg_out[7] ),
    .A1(\alu_out_q[7] ),
    .S(latched_stalu),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _41589_ (.A0(\reg_next_pc[6] ),
    .A1(_01479_),
    .S(latched_store),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _41590_ (.A0(\reg_out[6] ),
    .A1(\alu_out_q[6] ),
    .S(latched_stalu),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _41591_ (.A0(\reg_next_pc[5] ),
    .A1(_01476_),
    .S(latched_store),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _41592_ (.A0(\reg_out[5] ),
    .A1(\alu_out_q[5] ),
    .S(latched_stalu),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_2 _41593_ (.A0(_01474_),
    .A1(_01471_),
    .S(_00292_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _41594_ (.A0(\reg_next_pc[4] ),
    .A1(_01472_),
    .S(latched_store),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _41595_ (.A0(\reg_out[4] ),
    .A1(\alu_out_q[4] ),
    .S(latched_stalu),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _41596_ (.A0(\reg_next_pc[3] ),
    .A1(_01468_),
    .S(latched_store),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _41597_ (.A0(\reg_out[3] ),
    .A1(\alu_out_q[3] ),
    .S(latched_stalu),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _41598_ (.A0(\reg_next_pc[1] ),
    .A1(_01465_),
    .S(latched_store),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_2 _41599_ (.A0(\reg_out[1] ),
    .A1(\alu_out_q[1] ),
    .S(latched_stalu),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _41600_ (.A0(_01301_),
    .A1(\timer[31] ),
    .S(_01208_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _41601_ (.A0(_01298_),
    .A1(\timer[30] ),
    .S(_01208_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _41602_ (.A0(_01295_),
    .A1(\timer[29] ),
    .S(_01208_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _41603_ (.A0(_01292_),
    .A1(\timer[28] ),
    .S(_01208_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _41604_ (.A0(_01289_),
    .A1(\timer[27] ),
    .S(_01208_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _41605_ (.A0(_01286_),
    .A1(\timer[26] ),
    .S(_01208_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _41606_ (.A0(_01283_),
    .A1(\timer[25] ),
    .S(_01208_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _41607_ (.A0(_01280_),
    .A1(\timer[24] ),
    .S(_01208_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _41608_ (.A0(_01277_),
    .A1(\timer[23] ),
    .S(_01208_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _41609_ (.A0(_01274_),
    .A1(\timer[22] ),
    .S(_01208_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _41610_ (.A0(_01271_),
    .A1(\timer[21] ),
    .S(_01208_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _41611_ (.A0(_01268_),
    .A1(\timer[20] ),
    .S(_01208_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _41612_ (.A0(_01265_),
    .A1(\timer[19] ),
    .S(_01208_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _41613_ (.A0(_01262_),
    .A1(\timer[18] ),
    .S(_01208_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _41614_ (.A0(_01259_),
    .A1(\timer[17] ),
    .S(_01208_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _41615_ (.A0(_01256_),
    .A1(\timer[16] ),
    .S(_01208_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _41616_ (.A0(_01253_),
    .A1(\timer[15] ),
    .S(_01208_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _41617_ (.A0(_01250_),
    .A1(\timer[14] ),
    .S(_01208_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _41618_ (.A0(_01247_),
    .A1(\timer[13] ),
    .S(_01208_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _41619_ (.A0(_01244_),
    .A1(\timer[12] ),
    .S(_01208_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _41620_ (.A0(_01241_),
    .A1(\timer[11] ),
    .S(_01208_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _41621_ (.A0(_01238_),
    .A1(\timer[10] ),
    .S(_01208_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _41622_ (.A0(_01235_),
    .A1(\timer[9] ),
    .S(_01208_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _41623_ (.A0(_01232_),
    .A1(\timer[8] ),
    .S(_01208_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _41624_ (.A0(_01229_),
    .A1(\timer[7] ),
    .S(_01208_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _41625_ (.A0(_01226_),
    .A1(\timer[6] ),
    .S(_01208_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _41626_ (.A0(_01223_),
    .A1(\timer[5] ),
    .S(_01208_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _41627_ (.A0(_01220_),
    .A1(\timer[4] ),
    .S(_01208_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _41628_ (.A0(_01217_),
    .A1(\timer[3] ),
    .S(_01208_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _41629_ (.A0(_01214_),
    .A1(\timer[2] ),
    .S(_01208_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _41630_ (.A0(_01211_),
    .A1(\timer[1] ),
    .S(_01208_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_2 _41631_ (.A0(_01206_),
    .A1(_01201_),
    .S(net467),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_4 _41632_ (.A0(_01179_),
    .A1(_01174_),
    .S(net467),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_2 _41633_ (.A0(_01152_),
    .A1(_01147_),
    .S(net467),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_4 _41634_ (.A0(_01125_),
    .A1(_01120_),
    .S(net467),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_4 _41635_ (.A0(_01098_),
    .A1(_01093_),
    .S(net467),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_2 _41636_ (.A0(_01071_),
    .A1(_01066_),
    .S(net467),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_4 _41637_ (.A0(_01044_),
    .A1(_01039_),
    .S(net467),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_4 _41638_ (.A0(_01017_),
    .A1(_01012_),
    .S(net467),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_4 _41639_ (.A0(_00990_),
    .A1(_00985_),
    .S(net467),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_4 _41640_ (.A0(_00963_),
    .A1(_00958_),
    .S(net467),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_4 _41641_ (.A0(_00936_),
    .A1(_00931_),
    .S(net467),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_4 _41642_ (.A0(_00909_),
    .A1(_00904_),
    .S(net467),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_8 _41643_ (.A0(_00882_),
    .A1(_00877_),
    .S(_00368_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_8 _41644_ (.A0(_00855_),
    .A1(_00850_),
    .S(_00368_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_4 _41645_ (.A0(_00828_),
    .A1(_00823_),
    .S(_00368_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_8 _41646_ (.A0(_00801_),
    .A1(_00796_),
    .S(_00368_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_4 _41647_ (.A0(_00774_),
    .A1(_00769_),
    .S(_00368_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_4 _41648_ (.A0(_00747_),
    .A1(_00742_),
    .S(_00368_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_4 _41649_ (.A0(_00720_),
    .A1(_00715_),
    .S(net466),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_4 _41650_ (.A0(_00693_),
    .A1(_00688_),
    .S(net466),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_8 _41651_ (.A0(_00666_),
    .A1(_00661_),
    .S(net466),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_8 _41652_ (.A0(_00639_),
    .A1(_00634_),
    .S(net466),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_4 _41653_ (.A0(_00612_),
    .A1(_00607_),
    .S(net466),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_4 _41654_ (.A0(_00585_),
    .A1(_00580_),
    .S(net466),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_4 _41655_ (.A0(_00558_),
    .A1(_00553_),
    .S(net466),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_8 _41656_ (.A0(_00531_),
    .A1(_00526_),
    .S(net466),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_4 _41657_ (.A0(_00504_),
    .A1(_00499_),
    .S(net466),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_8 _41658_ (.A0(_00477_),
    .A1(_00472_),
    .S(net466),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_4 _41659_ (.A0(_00450_),
    .A1(_00445_),
    .S(net466),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_4 _41660_ (.A0(_00423_),
    .A1(_00418_),
    .S(net466),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_4 _41661_ (.A0(_00396_),
    .A1(_00391_),
    .S(_00368_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_2 _41662_ (.A0(_00369_),
    .A1(_00365_),
    .S(net467),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_8 _41663_ (.A0(_00366_),
    .A1(_00367_),
    .S(net507),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_8 _41664_ (.A0(\decoded_rs1[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(\cpu_state[3] ),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_4 _41665_ (.A0(\decoded_rs1[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(\cpu_state[3] ),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_4 _41666_ (.A0(\decoded_rs1[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(\cpu_state[3] ),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_8 _41667_ (.A0(\decoded_rs1[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(\cpu_state[3] ),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _41668_ (.A0(_00349_),
    .A1(_00323_),
    .S(decoder_trigger),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _41669_ (.A0(_00350_),
    .A1(_00351_),
    .S(_00309_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _41670_ (.A0(_00352_),
    .A1(_00349_),
    .S(_00308_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _41671_ (.A0(_00355_),
    .A1(_00353_),
    .S(_00354_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _41672_ (.A0(_00337_),
    .A1(_00344_),
    .S(is_beq_bne_blt_bge_bltu_bgeu),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _41673_ (.A0(_00345_),
    .A1(_00337_),
    .S(alu_wait),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_4 _41674_ (.A0(_00342_),
    .A1(_00340_),
    .S(_00341_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _41675_ (.A0(_00338_),
    .A1(_00337_),
    .S(_00296_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _41676_ (.A0(\mem_rdata_q[12] ),
    .A1(_00334_),
    .S(\mem_rdata_q[13] ),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _41677_ (.A0(\cpu_state[1] ),
    .A1(_00302_),
    .S(\cpu_state[4] ),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _41678_ (.A0(_00322_),
    .A1(_00296_),
    .S(\cpu_state[6] ),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _41679_ (.A0(_00315_),
    .A1(alu_wait),
    .S(\cpu_state[4] ),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _41680_ (.A0(\mem_rdata_q[6] ),
    .A1(net61),
    .S(mem_xfer),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_2 _41681_ (.A0(\mem_rdata_q[5] ),
    .A1(net512),
    .S(mem_xfer),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_2 _41682_ (.A0(\mem_rdata_q[4] ),
    .A1(net59),
    .S(mem_xfer),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _41683_ (.A0(\mem_rdata_q[3] ),
    .A1(net58),
    .S(mem_xfer),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _41684_ (.A0(\mem_rdata_q[2] ),
    .A1(net55),
    .S(net479),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _41685_ (.A0(\mem_rdata_q[1] ),
    .A1(net44),
    .S(net479),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _41686_ (.A0(\mem_rdata_q[0] ),
    .A1(net33),
    .S(net479),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _41687_ (.A0(\cpu_state[1] ),
    .A1(instr_retirq),
    .S(net508),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _41688_ (.A0(_00319_),
    .A1(\cpu_state[5] ),
    .S(_00296_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _41689_ (.A0(_00317_),
    .A1(\cpu_state[6] ),
    .S(_00296_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _41690_ (.A0(_00313_),
    .A1(_00312_),
    .S(_00307_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _41691_ (.A0(_00298_),
    .A1(_00299_),
    .S(_00289_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _41692_ (.A0(\reg_next_pc[2] ),
    .A1(_00293_),
    .S(latched_store),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _41693_ (.A0(\reg_out[2] ),
    .A1(\alu_out_q[2] ),
    .S(latched_stalu),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _41694_ (.A0(_00126_),
    .A1(_00122_),
    .S(net503),
    .X(_02558_));
 sky130_fd_sc_hd__mux2_1 _41695_ (.A0(_00120_),
    .A1(_00116_),
    .S(net225),
    .X(_02557_));
 sky130_fd_sc_hd__mux2_1 _41696_ (.A0(_00114_),
    .A1(_00110_),
    .S(net503),
    .X(_02556_));
 sky130_fd_sc_hd__mux2_1 _41697_ (.A0(_00108_),
    .A1(_00104_),
    .S(net225),
    .X(_02555_));
 sky130_fd_sc_hd__mux2_1 _41698_ (.A0(_00102_),
    .A1(_00095_),
    .S(net503),
    .X(_02554_));
 sky130_fd_sc_hd__mux2_1 _41699_ (.A0(_00092_),
    .A1(_00085_),
    .S(net503),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _41700_ (.A0(_00082_),
    .A1(_00068_),
    .S(net503),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _41701_ (.A0(_00064_),
    .A1(_00050_),
    .S(net225),
    .X(_02551_));
 sky130_fd_sc_hd__mux2_1 _41702_ (.A0(_01694_),
    .A1(_01695_),
    .S(_00290_),
    .X(_02541_));
 sky130_fd_sc_hd__mux2_1 _41703_ (.A0(_01691_),
    .A1(_01692_),
    .S(_00290_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _41704_ (.A0(_01688_),
    .A1(_01689_),
    .S(_00290_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _41705_ (.A0(_01685_),
    .A1(_01686_),
    .S(_00290_),
    .X(_02538_));
 sky130_fd_sc_hd__mux2_1 _41706_ (.A0(_01679_),
    .A1(_01680_),
    .S(instr_jal),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _41707_ (.A0(_01682_),
    .A1(_02581_),
    .S(net412),
    .X(_02530_));
 sky130_fd_sc_hd__mux2_1 _41708_ (.A0(_01675_),
    .A1(_01676_),
    .S(instr_jal),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _41709_ (.A0(_01678_),
    .A1(_02580_),
    .S(net412),
    .X(_02529_));
 sky130_fd_sc_hd__mux2_1 _41710_ (.A0(_01671_),
    .A1(_01672_),
    .S(instr_jal),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _41711_ (.A0(_01674_),
    .A1(_02579_),
    .S(net412),
    .X(_02527_));
 sky130_fd_sc_hd__mux2_1 _41712_ (.A0(_01667_),
    .A1(_01668_),
    .S(instr_jal),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _41713_ (.A0(_01670_),
    .A1(_02578_),
    .S(net412),
    .X(_02526_));
 sky130_fd_sc_hd__mux2_1 _41714_ (.A0(_01663_),
    .A1(_01664_),
    .S(instr_jal),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _41715_ (.A0(_01666_),
    .A1(_02577_),
    .S(net412),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _41716_ (.A0(_01659_),
    .A1(_01660_),
    .S(instr_jal),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _41717_ (.A0(_01662_),
    .A1(_02576_),
    .S(net412),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _41718_ (.A0(_01655_),
    .A1(_01656_),
    .S(instr_jal),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _41719_ (.A0(_01658_),
    .A1(_02575_),
    .S(net412),
    .X(_02523_));
 sky130_fd_sc_hd__mux2_1 _41720_ (.A0(_01651_),
    .A1(_01652_),
    .S(instr_jal),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _41721_ (.A0(_01654_),
    .A1(_02574_),
    .S(net412),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _41722_ (.A0(_01647_),
    .A1(_01648_),
    .S(instr_jal),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _41723_ (.A0(_01650_),
    .A1(_02573_),
    .S(net412),
    .X(_02521_));
 sky130_fd_sc_hd__mux2_1 _41724_ (.A0(_01643_),
    .A1(_01644_),
    .S(instr_jal),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _41725_ (.A0(_01646_),
    .A1(_02572_),
    .S(net412),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _41726_ (.A0(_01639_),
    .A1(_01640_),
    .S(instr_jal),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _41727_ (.A0(_01642_),
    .A1(_02570_),
    .S(net412),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _41728_ (.A0(_01635_),
    .A1(_01636_),
    .S(instr_jal),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _41729_ (.A0(_01638_),
    .A1(_02569_),
    .S(net412),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _41730_ (.A0(_01631_),
    .A1(_01632_),
    .S(instr_jal),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _41731_ (.A0(_01634_),
    .A1(_02568_),
    .S(net412),
    .X(_02516_));
 sky130_fd_sc_hd__mux2_1 _41732_ (.A0(_01627_),
    .A1(_01628_),
    .S(instr_jal),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _41733_ (.A0(_01630_),
    .A1(_02567_),
    .S(net412),
    .X(_02515_));
 sky130_fd_sc_hd__mux2_1 _41734_ (.A0(_01623_),
    .A1(_01624_),
    .S(instr_jal),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _41735_ (.A0(_01626_),
    .A1(_02566_),
    .S(net412),
    .X(_02514_));
 sky130_fd_sc_hd__mux2_1 _41736_ (.A0(_01619_),
    .A1(_01620_),
    .S(instr_jal),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _41737_ (.A0(_01622_),
    .A1(_02565_),
    .S(net412),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _41738_ (.A0(_01615_),
    .A1(_01616_),
    .S(instr_jal),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _41739_ (.A0(_01618_),
    .A1(_02564_),
    .S(net412),
    .X(_02512_));
 sky130_fd_sc_hd__mux2_1 _41740_ (.A0(_01611_),
    .A1(_01612_),
    .S(instr_jal),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _41741_ (.A0(_01614_),
    .A1(_02563_),
    .S(net413),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _41742_ (.A0(_01607_),
    .A1(_01608_),
    .S(instr_jal),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _41743_ (.A0(_01610_),
    .A1(_02562_),
    .S(net413),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _41744_ (.A0(_01603_),
    .A1(_01604_),
    .S(instr_jal),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _41745_ (.A0(_01606_),
    .A1(_02561_),
    .S(net413),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _41746_ (.A0(_01599_),
    .A1(_01600_),
    .S(instr_jal),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _41747_ (.A0(_01602_),
    .A1(_02589_),
    .S(net413),
    .X(_02508_));
 sky130_fd_sc_hd__mux2_1 _41748_ (.A0(_01595_),
    .A1(_01596_),
    .S(instr_jal),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _41749_ (.A0(_01598_),
    .A1(_02588_),
    .S(net413),
    .X(_02507_));
 sky130_fd_sc_hd__mux2_1 _41750_ (.A0(_01591_),
    .A1(_01592_),
    .S(instr_jal),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _41751_ (.A0(_01594_),
    .A1(_02587_),
    .S(net413),
    .X(_02537_));
 sky130_fd_sc_hd__mux2_1 _41752_ (.A0(_01587_),
    .A1(_01588_),
    .S(instr_jal),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _41753_ (.A0(_01590_),
    .A1(_02586_),
    .S(net413),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _41754_ (.A0(_01583_),
    .A1(_01584_),
    .S(instr_jal),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _41755_ (.A0(_01586_),
    .A1(_02585_),
    .S(net413),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _41756_ (.A0(_01579_),
    .A1(_01580_),
    .S(instr_jal),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _41757_ (.A0(_01582_),
    .A1(_02584_),
    .S(net413),
    .X(_02534_));
 sky130_fd_sc_hd__mux2_1 _41758_ (.A0(_01575_),
    .A1(_01576_),
    .S(instr_jal),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _41759_ (.A0(_01578_),
    .A1(_02583_),
    .S(net413),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _41760_ (.A0(_01571_),
    .A1(_01572_),
    .S(instr_jal),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _41761_ (.A0(_01574_),
    .A1(_02582_),
    .S(net413),
    .X(_02532_));
 sky130_fd_sc_hd__mux2_1 _41762_ (.A0(_01567_),
    .A1(_01568_),
    .S(instr_jal),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _41763_ (.A0(_01570_),
    .A1(_02571_),
    .S(net413),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _41764_ (.A0(_01561_),
    .A1(_01562_),
    .S(instr_jal),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _41765_ (.A0(_02560_),
    .A1(_01563_),
    .S(decoder_trigger),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _41766_ (.A0(_01564_),
    .A1(_01565_),
    .S(_00309_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _41767_ (.A0(_01566_),
    .A1(_02560_),
    .S(net413),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _41768_ (.A0(_02590_),
    .A1(_01557_),
    .S(instr_jal),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _41769_ (.A0(_02590_),
    .A1(_01558_),
    .S(decoder_trigger),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _41770_ (.A0(_01559_),
    .A1(_02590_),
    .S(_00309_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _41771_ (.A0(_01560_),
    .A1(_02590_),
    .S(net413),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_2 _41772_ (.A0(\cpuregs_rs1[31] ),
    .A1(_01462_),
    .S(is_lui_auipc_jal),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _41773_ (.A0(_01464_),
    .A1(_01463_),
    .S(net501),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _41774_ (.A0(\cpuregs_rs1[30] ),
    .A1(_01459_),
    .S(is_lui_auipc_jal),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _41775_ (.A0(_01461_),
    .A1(_01460_),
    .S(net501),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _41776_ (.A0(\cpuregs_rs1[29] ),
    .A1(_01456_),
    .S(is_lui_auipc_jal),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _41777_ (.A0(_01458_),
    .A1(_01457_),
    .S(net501),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _41778_ (.A0(\cpuregs_rs1[28] ),
    .A1(_01453_),
    .S(is_lui_auipc_jal),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _41779_ (.A0(_01455_),
    .A1(_01454_),
    .S(net501),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _41780_ (.A0(\cpuregs_rs1[27] ),
    .A1(_01450_),
    .S(is_lui_auipc_jal),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _41781_ (.A0(_01452_),
    .A1(_01451_),
    .S(net501),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _41782_ (.A0(\cpuregs_rs1[26] ),
    .A1(_01447_),
    .S(is_lui_auipc_jal),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _41783_ (.A0(_01449_),
    .A1(_01448_),
    .S(net501),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _41784_ (.A0(\cpuregs_rs1[25] ),
    .A1(_01444_),
    .S(is_lui_auipc_jal),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _41785_ (.A0(_01446_),
    .A1(_01445_),
    .S(net501),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _41786_ (.A0(\cpuregs_rs1[24] ),
    .A1(_01441_),
    .S(is_lui_auipc_jal),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _41787_ (.A0(_01443_),
    .A1(_01442_),
    .S(net501),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _41788_ (.A0(\cpuregs_rs1[23] ),
    .A1(_01438_),
    .S(is_lui_auipc_jal),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _41789_ (.A0(_01440_),
    .A1(_01439_),
    .S(net501),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _41790_ (.A0(\cpuregs_rs1[22] ),
    .A1(_01435_),
    .S(is_lui_auipc_jal),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _41791_ (.A0(_01437_),
    .A1(_01436_),
    .S(net500),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _41792_ (.A0(\cpuregs_rs1[21] ),
    .A1(_01432_),
    .S(is_lui_auipc_jal),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _41793_ (.A0(_01434_),
    .A1(_01433_),
    .S(net500),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _41794_ (.A0(\cpuregs_rs1[20] ),
    .A1(_01429_),
    .S(is_lui_auipc_jal),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _41795_ (.A0(_01431_),
    .A1(_01430_),
    .S(net500),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _41796_ (.A0(\cpuregs_rs1[19] ),
    .A1(_01426_),
    .S(is_lui_auipc_jal),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _41797_ (.A0(_01428_),
    .A1(_01427_),
    .S(net500),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _41798_ (.A0(\cpuregs_rs1[18] ),
    .A1(_01423_),
    .S(is_lui_auipc_jal),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _41799_ (.A0(_01425_),
    .A1(_01424_),
    .S(net500),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _41800_ (.A0(\cpuregs_rs1[17] ),
    .A1(_01420_),
    .S(is_lui_auipc_jal),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _41801_ (.A0(_01422_),
    .A1(_01421_),
    .S(net500),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _41802_ (.A0(\cpuregs_rs1[16] ),
    .A1(_01417_),
    .S(is_lui_auipc_jal),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _41803_ (.A0(_01419_),
    .A1(_01418_),
    .S(net500),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _41804_ (.A0(\cpuregs_rs1[15] ),
    .A1(_01414_),
    .S(is_lui_auipc_jal),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _41805_ (.A0(_01416_),
    .A1(_01415_),
    .S(net500),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _41806_ (.A0(\cpuregs_rs1[14] ),
    .A1(_01411_),
    .S(is_lui_auipc_jal),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _41807_ (.A0(_01413_),
    .A1(_01412_),
    .S(net500),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _41808_ (.A0(\cpuregs_rs1[13] ),
    .A1(_01408_),
    .S(is_lui_auipc_jal),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _41809_ (.A0(_01410_),
    .A1(_01409_),
    .S(net500),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _41810_ (.A0(\cpuregs_rs1[12] ),
    .A1(_01405_),
    .S(is_lui_auipc_jal),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _41811_ (.A0(_01407_),
    .A1(_01406_),
    .S(net500),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _41812_ (.A0(\cpuregs_rs1[11] ),
    .A1(_01402_),
    .S(is_lui_auipc_jal),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _41813_ (.A0(_01404_),
    .A1(_01403_),
    .S(net500),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _41814_ (.A0(\cpuregs_rs1[10] ),
    .A1(_01399_),
    .S(is_lui_auipc_jal),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _41815_ (.A0(_01401_),
    .A1(_01400_),
    .S(net500),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _41816_ (.A0(\cpuregs_rs1[9] ),
    .A1(_01396_),
    .S(is_lui_auipc_jal),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _41817_ (.A0(_01398_),
    .A1(_01397_),
    .S(net500),
    .X(_02506_));
 sky130_fd_sc_hd__mux2_1 _41818_ (.A0(\cpuregs_rs1[8] ),
    .A1(_01393_),
    .S(is_lui_auipc_jal),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _41819_ (.A0(_01395_),
    .A1(_01394_),
    .S(net500),
    .X(_02505_));
 sky130_fd_sc_hd__mux2_1 _41820_ (.A0(\cpuregs_rs1[7] ),
    .A1(_01390_),
    .S(is_lui_auipc_jal),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _41821_ (.A0(_01392_),
    .A1(_01391_),
    .S(net500),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _41822_ (.A0(\cpuregs_rs1[6] ),
    .A1(_01387_),
    .S(is_lui_auipc_jal),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _41823_ (.A0(_01389_),
    .A1(_01388_),
    .S(net500),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_1 _41824_ (.A0(\cpuregs_rs1[5] ),
    .A1(_01384_),
    .S(is_lui_auipc_jal),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _41825_ (.A0(_01386_),
    .A1(_01385_),
    .S(net500),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _41826_ (.A0(\cpuregs_rs1[4] ),
    .A1(_01381_),
    .S(is_lui_auipc_jal),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _41827_ (.A0(_01383_),
    .A1(_01382_),
    .S(net501),
    .X(_02501_));
 sky130_fd_sc_hd__mux2_1 _41828_ (.A0(\cpuregs_rs1[3] ),
    .A1(_01378_),
    .S(is_lui_auipc_jal),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _41829_ (.A0(_01380_),
    .A1(_01379_),
    .S(net501),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _41830_ (.A0(\cpuregs_rs1[2] ),
    .A1(_01375_),
    .S(is_lui_auipc_jal),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _41831_ (.A0(_01377_),
    .A1(_01376_),
    .S(net501),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _41832_ (.A0(\cpuregs_rs1[1] ),
    .A1(_01372_),
    .S(is_lui_auipc_jal),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _41833_ (.A0(_01374_),
    .A1(_01373_),
    .S(net501),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _41834_ (.A0(\cpuregs_rs1[0] ),
    .A1(_01369_),
    .S(is_lui_auipc_jal),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _41835_ (.A0(_01371_),
    .A1(_01370_),
    .S(net501),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _41836_ (.A0(_01367_),
    .A1(\decoded_imm[31] ),
    .S(_01304_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _41837_ (.A0(_01368_),
    .A1(\cpuregs_rs1[31] ),
    .S(net507),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _41838_ (.A0(_01365_),
    .A1(\decoded_imm[30] ),
    .S(_01304_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _41839_ (.A0(_01366_),
    .A1(\cpuregs_rs1[30] ),
    .S(\cpu_state[3] ),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _41840_ (.A0(_01363_),
    .A1(\decoded_imm[29] ),
    .S(_01304_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _41841_ (.A0(_01364_),
    .A1(\cpuregs_rs1[29] ),
    .S(\cpu_state[3] ),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _41842_ (.A0(_01361_),
    .A1(\decoded_imm[28] ),
    .S(_01304_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _41843_ (.A0(_01362_),
    .A1(\cpuregs_rs1[28] ),
    .S(net507),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _41844_ (.A0(_01359_),
    .A1(\decoded_imm[27] ),
    .S(_01304_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _41845_ (.A0(_01360_),
    .A1(\cpuregs_rs1[27] ),
    .S(net507),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _41846_ (.A0(_01357_),
    .A1(\decoded_imm[26] ),
    .S(_01304_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _41847_ (.A0(_01358_),
    .A1(\cpuregs_rs1[26] ),
    .S(net507),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _41848_ (.A0(_01355_),
    .A1(\decoded_imm[25] ),
    .S(_01304_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _41849_ (.A0(_01356_),
    .A1(\cpuregs_rs1[25] ),
    .S(net507),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _41850_ (.A0(_01353_),
    .A1(\decoded_imm[24] ),
    .S(_01304_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _41851_ (.A0(_01354_),
    .A1(\cpuregs_rs1[24] ),
    .S(net507),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _41852_ (.A0(_01351_),
    .A1(\decoded_imm[23] ),
    .S(net475),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _41853_ (.A0(_01352_),
    .A1(\cpuregs_rs1[23] ),
    .S(net507),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _41854_ (.A0(_01349_),
    .A1(\decoded_imm[22] ),
    .S(net475),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _41855_ (.A0(_01350_),
    .A1(\cpuregs_rs1[22] ),
    .S(net507),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _41856_ (.A0(_01347_),
    .A1(\decoded_imm[21] ),
    .S(net475),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _41857_ (.A0(_01348_),
    .A1(\cpuregs_rs1[21] ),
    .S(net507),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _41858_ (.A0(_01345_),
    .A1(\decoded_imm[20] ),
    .S(net475),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _41859_ (.A0(_01346_),
    .A1(\cpuregs_rs1[20] ),
    .S(net507),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _41860_ (.A0(_01343_),
    .A1(\decoded_imm[19] ),
    .S(net475),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _41861_ (.A0(_01344_),
    .A1(\cpuregs_rs1[19] ),
    .S(net507),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _41862_ (.A0(_01341_),
    .A1(\decoded_imm[18] ),
    .S(net475),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _41863_ (.A0(_01342_),
    .A1(\cpuregs_rs1[18] ),
    .S(net507),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _41864_ (.A0(_01339_),
    .A1(\decoded_imm[17] ),
    .S(net475),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _41865_ (.A0(_01340_),
    .A1(\cpuregs_rs1[17] ),
    .S(net507),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _41866_ (.A0(_01337_),
    .A1(\decoded_imm[16] ),
    .S(net475),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _41867_ (.A0(_01338_),
    .A1(\cpuregs_rs1[16] ),
    .S(net507),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _41868_ (.A0(_01335_),
    .A1(\decoded_imm[15] ),
    .S(net475),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _41869_ (.A0(_01336_),
    .A1(\cpuregs_rs1[15] ),
    .S(net507),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _41870_ (.A0(_01333_),
    .A1(\decoded_imm[14] ),
    .S(net475),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _41871_ (.A0(_01334_),
    .A1(\cpuregs_rs1[14] ),
    .S(net507),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _41872_ (.A0(_01331_),
    .A1(\decoded_imm[13] ),
    .S(net475),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _41873_ (.A0(_01332_),
    .A1(\cpuregs_rs1[13] ),
    .S(net507),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _41874_ (.A0(_01329_),
    .A1(\decoded_imm[12] ),
    .S(net475),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _41875_ (.A0(_01330_),
    .A1(\cpuregs_rs1[12] ),
    .S(net507),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _41876_ (.A0(_01327_),
    .A1(\decoded_imm[11] ),
    .S(net475),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _41877_ (.A0(_01328_),
    .A1(\cpuregs_rs1[11] ),
    .S(net507),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _41878_ (.A0(_01325_),
    .A1(\decoded_imm[10] ),
    .S(net475),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _41879_ (.A0(_01326_),
    .A1(\cpuregs_rs1[10] ),
    .S(net507),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _41880_ (.A0(_01323_),
    .A1(\decoded_imm[9] ),
    .S(net475),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _41881_ (.A0(_01324_),
    .A1(\cpuregs_rs1[9] ),
    .S(net507),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _41882_ (.A0(_01321_),
    .A1(\decoded_imm[8] ),
    .S(net475),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _41883_ (.A0(_01322_),
    .A1(\cpuregs_rs1[8] ),
    .S(net507),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _41884_ (.A0(_01319_),
    .A1(\decoded_imm[7] ),
    .S(net475),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _41885_ (.A0(_01320_),
    .A1(\cpuregs_rs1[7] ),
    .S(net507),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _41886_ (.A0(_01317_),
    .A1(\decoded_imm[6] ),
    .S(net475),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _41887_ (.A0(_01318_),
    .A1(\cpuregs_rs1[6] ),
    .S(net507),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _41888_ (.A0(_01315_),
    .A1(\decoded_imm[5] ),
    .S(net475),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _41889_ (.A0(_01316_),
    .A1(\cpuregs_rs1[5] ),
    .S(net507),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _41890_ (.A0(\decoded_imm[4] ),
    .A1(\decoded_imm_uj[4] ),
    .S(is_slli_srli_srai),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _41891_ (.A0(_01313_),
    .A1(\decoded_imm[4] ),
    .S(_01304_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _41892_ (.A0(_01314_),
    .A1(\cpuregs_rs1[4] ),
    .S(net507),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _41893_ (.A0(\decoded_imm[3] ),
    .A1(\decoded_imm_uj[3] ),
    .S(is_slli_srli_srai),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _41894_ (.A0(_01311_),
    .A1(\decoded_imm[3] ),
    .S(_01304_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _41895_ (.A0(_01312_),
    .A1(\cpuregs_rs1[3] ),
    .S(net507),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _41896_ (.A0(\decoded_imm[2] ),
    .A1(\decoded_imm_uj[2] ),
    .S(is_slli_srli_srai),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _41897_ (.A0(_01309_),
    .A1(\decoded_imm[2] ),
    .S(_01304_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _41898_ (.A0(_01310_),
    .A1(\cpuregs_rs1[2] ),
    .S(net507),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _41899_ (.A0(\decoded_imm[1] ),
    .A1(\decoded_imm_uj[1] ),
    .S(is_slli_srli_srai),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _41900_ (.A0(_01307_),
    .A1(\decoded_imm[1] ),
    .S(_01304_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _41901_ (.A0(_01308_),
    .A1(\cpuregs_rs1[1] ),
    .S(net507),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _41902_ (.A0(\decoded_imm[0] ),
    .A1(\decoded_imm_uj[11] ),
    .S(is_slli_srli_srai),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _41903_ (.A0(_01305_),
    .A1(\decoded_imm[0] ),
    .S(_01304_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _41904_ (.A0(_01306_),
    .A1(\cpuregs_rs1[0] ),
    .S(net507),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _41905_ (.A0(_01302_),
    .A1(\cpuregs_rs1[31] ),
    .S(instr_timer),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _41906_ (.A0(_01302_),
    .A1(_01303_),
    .S(\cpu_state[2] ),
    .X(_02435_));
 sky130_fd_sc_hd__mux2_1 _41907_ (.A0(_01299_),
    .A1(\cpuregs_rs1[30] ),
    .S(instr_timer),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _41908_ (.A0(_01299_),
    .A1(_01300_),
    .S(\cpu_state[2] ),
    .X(_02434_));
 sky130_fd_sc_hd__mux2_1 _41909_ (.A0(_01296_),
    .A1(\cpuregs_rs1[29] ),
    .S(instr_timer),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _41910_ (.A0(_01296_),
    .A1(_01297_),
    .S(\cpu_state[2] ),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _41911_ (.A0(_01293_),
    .A1(\cpuregs_rs1[28] ),
    .S(instr_timer),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _41912_ (.A0(_01293_),
    .A1(_01294_),
    .S(\cpu_state[2] ),
    .X(_02431_));
 sky130_fd_sc_hd__mux2_1 _41913_ (.A0(_01290_),
    .A1(\cpuregs_rs1[27] ),
    .S(instr_timer),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _41914_ (.A0(_01290_),
    .A1(_01291_),
    .S(\cpu_state[2] ),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _41915_ (.A0(_01287_),
    .A1(\cpuregs_rs1[26] ),
    .S(instr_timer),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _41916_ (.A0(_01287_),
    .A1(_01288_),
    .S(\cpu_state[2] ),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _41917_ (.A0(_01284_),
    .A1(\cpuregs_rs1[25] ),
    .S(instr_timer),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _41918_ (.A0(_01284_),
    .A1(_01285_),
    .S(\cpu_state[2] ),
    .X(_02428_));
 sky130_fd_sc_hd__mux2_1 _41919_ (.A0(_01281_),
    .A1(\cpuregs_rs1[24] ),
    .S(instr_timer),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _41920_ (.A0(_01281_),
    .A1(_01282_),
    .S(\cpu_state[2] ),
    .X(_02427_));
 sky130_fd_sc_hd__mux2_1 _41921_ (.A0(_01278_),
    .A1(\cpuregs_rs1[23] ),
    .S(instr_timer),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _41922_ (.A0(_01278_),
    .A1(_01279_),
    .S(\cpu_state[2] ),
    .X(_02426_));
 sky130_fd_sc_hd__mux2_1 _41923_ (.A0(_01275_),
    .A1(\cpuregs_rs1[22] ),
    .S(instr_timer),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _41924_ (.A0(_01275_),
    .A1(_01276_),
    .S(\cpu_state[2] ),
    .X(_02425_));
 sky130_fd_sc_hd__mux2_1 _41925_ (.A0(_01272_),
    .A1(\cpuregs_rs1[21] ),
    .S(instr_timer),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _41926_ (.A0(_01272_),
    .A1(_01273_),
    .S(\cpu_state[2] ),
    .X(_02424_));
 sky130_fd_sc_hd__mux2_1 _41927_ (.A0(_01269_),
    .A1(\cpuregs_rs1[20] ),
    .S(instr_timer),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _41928_ (.A0(_01269_),
    .A1(_01270_),
    .S(\cpu_state[2] ),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _41929_ (.A0(_01266_),
    .A1(\cpuregs_rs1[19] ),
    .S(instr_timer),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _41930_ (.A0(_01266_),
    .A1(_01267_),
    .S(\cpu_state[2] ),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _41931_ (.A0(_01263_),
    .A1(\cpuregs_rs1[18] ),
    .S(instr_timer),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _41932_ (.A0(_01263_),
    .A1(_01264_),
    .S(\cpu_state[2] ),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_1 _41933_ (.A0(_01260_),
    .A1(\cpuregs_rs1[17] ),
    .S(instr_timer),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _41934_ (.A0(_01260_),
    .A1(_01261_),
    .S(\cpu_state[2] ),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _41935_ (.A0(_01257_),
    .A1(\cpuregs_rs1[16] ),
    .S(instr_timer),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _41936_ (.A0(_01257_),
    .A1(_01258_),
    .S(\cpu_state[2] ),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _41937_ (.A0(_01254_),
    .A1(\cpuregs_rs1[15] ),
    .S(instr_timer),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _41938_ (.A0(_01254_),
    .A1(_01255_),
    .S(\cpu_state[2] ),
    .X(_02417_));
 sky130_fd_sc_hd__mux2_1 _41939_ (.A0(_01251_),
    .A1(\cpuregs_rs1[14] ),
    .S(instr_timer),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _41940_ (.A0(_01251_),
    .A1(_01252_),
    .S(\cpu_state[2] ),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _41941_ (.A0(_01248_),
    .A1(\cpuregs_rs1[13] ),
    .S(instr_timer),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _41942_ (.A0(_01248_),
    .A1(_01249_),
    .S(\cpu_state[2] ),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _41943_ (.A0(_01245_),
    .A1(\cpuregs_rs1[12] ),
    .S(instr_timer),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _41944_ (.A0(_01245_),
    .A1(_01246_),
    .S(\cpu_state[2] ),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _41945_ (.A0(_01242_),
    .A1(\cpuregs_rs1[11] ),
    .S(instr_timer),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _41946_ (.A0(_01242_),
    .A1(_01243_),
    .S(\cpu_state[2] ),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _41947_ (.A0(_01239_),
    .A1(\cpuregs_rs1[10] ),
    .S(instr_timer),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _41948_ (.A0(_01239_),
    .A1(_01240_),
    .S(net508),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _41949_ (.A0(_01236_),
    .A1(\cpuregs_rs1[9] ),
    .S(instr_timer),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _41950_ (.A0(_01236_),
    .A1(_01237_),
    .S(net508),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _41951_ (.A0(_01233_),
    .A1(\cpuregs_rs1[8] ),
    .S(instr_timer),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _41952_ (.A0(_01233_),
    .A1(_01234_),
    .S(net508),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _41953_ (.A0(_01230_),
    .A1(\cpuregs_rs1[7] ),
    .S(instr_timer),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _41954_ (.A0(_01230_),
    .A1(_01231_),
    .S(net508),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _41955_ (.A0(_01227_),
    .A1(\cpuregs_rs1[6] ),
    .S(instr_timer),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _41956_ (.A0(_01227_),
    .A1(_01228_),
    .S(net508),
    .X(_02439_));
 sky130_fd_sc_hd__mux2_1 _41957_ (.A0(_01224_),
    .A1(\cpuregs_rs1[5] ),
    .S(instr_timer),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _41958_ (.A0(_01224_),
    .A1(_01225_),
    .S(net508),
    .X(_02438_));
 sky130_fd_sc_hd__mux2_1 _41959_ (.A0(_01221_),
    .A1(\cpuregs_rs1[4] ),
    .S(instr_timer),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _41960_ (.A0(_01221_),
    .A1(_01222_),
    .S(net508),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _41961_ (.A0(_01218_),
    .A1(\cpuregs_rs1[3] ),
    .S(instr_timer),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _41962_ (.A0(_01218_),
    .A1(_01219_),
    .S(net508),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _41963_ (.A0(_01215_),
    .A1(\cpuregs_rs1[2] ),
    .S(instr_timer),
    .X(_01216_));
 sky130_fd_sc_hd__mux2_1 _41964_ (.A0(_01215_),
    .A1(_01216_),
    .S(net508),
    .X(_02433_));
 sky130_fd_sc_hd__mux2_1 _41965_ (.A0(_01212_),
    .A1(\cpuregs_rs1[1] ),
    .S(instr_timer),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _41966_ (.A0(_01212_),
    .A1(_01213_),
    .S(net508),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _41967_ (.A0(_01209_),
    .A1(\cpuregs_rs1[0] ),
    .S(instr_timer),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _41968_ (.A0(_01209_),
    .A1(_01210_),
    .S(net508),
    .X(_02411_));
 sky130_fd_sc_hd__mux4_1 _41969_ (.A0(_01202_),
    .A1(_01203_),
    .A2(_01204_),
    .A3(_01205_),
    .S0(_00357_),
    .S1(net482),
    .X(_01206_));
 sky130_fd_sc_hd__mux4_2 _41970_ (.A0(_01181_),
    .A1(_01182_),
    .A2(_01183_),
    .A3(_01184_),
    .S0(_00357_),
    .S1(net482),
    .X(_01185_));
 sky130_fd_sc_hd__mux4_1 _41971_ (.A0(_01186_),
    .A1(_01187_),
    .A2(_01188_),
    .A3(_01189_),
    .S0(_00357_),
    .S1(net482),
    .X(_01190_));
 sky130_fd_sc_hd__mux4_1 _41972_ (.A0(_01191_),
    .A1(_01192_),
    .A2(_01193_),
    .A3(_01194_),
    .S0(_00357_),
    .S1(net482),
    .X(_01195_));
 sky130_fd_sc_hd__mux4_1 _41973_ (.A0(_01196_),
    .A1(_01197_),
    .A2(_01198_),
    .A3(_01199_),
    .S0(_00357_),
    .S1(net482),
    .X(_01200_));
 sky130_fd_sc_hd__mux4_2 _41974_ (.A0(_01185_),
    .A1(_01190_),
    .A2(_01195_),
    .A3(_01200_),
    .S0(net490),
    .S1(net493),
    .X(_01201_));
 sky130_fd_sc_hd__mux4_1 _41975_ (.A0(_01175_),
    .A1(_01176_),
    .A2(_01177_),
    .A3(_01178_),
    .S0(_00357_),
    .S1(net481),
    .X(_01179_));
 sky130_fd_sc_hd__mux4_1 _41976_ (.A0(_01154_),
    .A1(_01155_),
    .A2(_01156_),
    .A3(_01157_),
    .S0(_00357_),
    .S1(net481),
    .X(_01158_));
 sky130_fd_sc_hd__mux4_2 _41977_ (.A0(_01159_),
    .A1(_01160_),
    .A2(_01161_),
    .A3(_01162_),
    .S0(_00357_),
    .S1(net481),
    .X(_01163_));
 sky130_fd_sc_hd__mux4_1 _41978_ (.A0(_01164_),
    .A1(_01165_),
    .A2(_01166_),
    .A3(_01167_),
    .S0(_00357_),
    .S1(net481),
    .X(_01168_));
 sky130_fd_sc_hd__mux4_2 _41979_ (.A0(_01169_),
    .A1(_01170_),
    .A2(_01171_),
    .A3(_01172_),
    .S0(_00357_),
    .S1(net481),
    .X(_01173_));
 sky130_fd_sc_hd__mux4_2 _41980_ (.A0(_01158_),
    .A1(_01163_),
    .A2(_01168_),
    .A3(_01173_),
    .S0(net490),
    .S1(_00362_),
    .X(_01174_));
 sky130_fd_sc_hd__mux4_1 _41981_ (.A0(_01148_),
    .A1(_01149_),
    .A2(_01150_),
    .A3(_01151_),
    .S0(_00357_),
    .S1(net481),
    .X(_01152_));
 sky130_fd_sc_hd__mux4_2 _41982_ (.A0(_01127_),
    .A1(_01128_),
    .A2(_01129_),
    .A3(_01130_),
    .S0(_00357_),
    .S1(net481),
    .X(_01131_));
 sky130_fd_sc_hd__mux4_1 _41983_ (.A0(_01132_),
    .A1(_01133_),
    .A2(_01134_),
    .A3(_01135_),
    .S0(_00357_),
    .S1(net481),
    .X(_01136_));
 sky130_fd_sc_hd__mux4_1 _41984_ (.A0(_01137_),
    .A1(_01138_),
    .A2(_01139_),
    .A3(_01140_),
    .S0(_00357_),
    .S1(net481),
    .X(_01141_));
 sky130_fd_sc_hd__mux4_2 _41985_ (.A0(_01142_),
    .A1(_01143_),
    .A2(_01144_),
    .A3(_01145_),
    .S0(_00357_),
    .S1(net481),
    .X(_01146_));
 sky130_fd_sc_hd__mux4_2 _41986_ (.A0(_01131_),
    .A1(_01136_),
    .A2(_01141_),
    .A3(_01146_),
    .S0(net490),
    .S1(net493),
    .X(_01147_));
 sky130_fd_sc_hd__mux4_2 _41987_ (.A0(_01121_),
    .A1(_01122_),
    .A2(_01123_),
    .A3(_01124_),
    .S0(_00357_),
    .S1(net481),
    .X(_01125_));
 sky130_fd_sc_hd__mux4_2 _41988_ (.A0(_01100_),
    .A1(_01101_),
    .A2(_01102_),
    .A3(_01103_),
    .S0(_00357_),
    .S1(net481),
    .X(_01104_));
 sky130_fd_sc_hd__mux4_1 _41989_ (.A0(_01105_),
    .A1(_01106_),
    .A2(_01107_),
    .A3(_01108_),
    .S0(_00357_),
    .S1(net481),
    .X(_01109_));
 sky130_fd_sc_hd__mux4_1 _41990_ (.A0(_01110_),
    .A1(_01111_),
    .A2(_01112_),
    .A3(_01113_),
    .S0(_00357_),
    .S1(net481),
    .X(_01114_));
 sky130_fd_sc_hd__mux4_2 _41991_ (.A0(_01115_),
    .A1(_01116_),
    .A2(_01117_),
    .A3(_01118_),
    .S0(_00357_),
    .S1(net481),
    .X(_01119_));
 sky130_fd_sc_hd__mux4_2 _41992_ (.A0(_01104_),
    .A1(_01109_),
    .A2(_01114_),
    .A3(_01119_),
    .S0(net490),
    .S1(_00362_),
    .X(_01120_));
 sky130_fd_sc_hd__mux4_1 _41993_ (.A0(_01094_),
    .A1(_01095_),
    .A2(_01096_),
    .A3(_01097_),
    .S0(_00357_),
    .S1(net481),
    .X(_01098_));
 sky130_fd_sc_hd__mux4_2 _41994_ (.A0(_01073_),
    .A1(_01074_),
    .A2(_01075_),
    .A3(_01076_),
    .S0(_00357_),
    .S1(net481),
    .X(_01077_));
 sky130_fd_sc_hd__mux4_1 _41995_ (.A0(_01078_),
    .A1(_01079_),
    .A2(_01080_),
    .A3(_01081_),
    .S0(_00357_),
    .S1(net481),
    .X(_01082_));
 sky130_fd_sc_hd__mux4_1 _41996_ (.A0(_01083_),
    .A1(_01084_),
    .A2(_01085_),
    .A3(_01086_),
    .S0(_00357_),
    .S1(net481),
    .X(_01087_));
 sky130_fd_sc_hd__mux4_2 _41997_ (.A0(_01088_),
    .A1(_01089_),
    .A2(_01090_),
    .A3(_01091_),
    .S0(_00357_),
    .S1(net481),
    .X(_01092_));
 sky130_fd_sc_hd__mux4_2 _41998_ (.A0(_01077_),
    .A1(_01082_),
    .A2(_01087_),
    .A3(_01092_),
    .S0(net490),
    .S1(_00362_),
    .X(_01093_));
 sky130_fd_sc_hd__mux4_1 _41999_ (.A0(_01067_),
    .A1(_01068_),
    .A2(_01069_),
    .A3(_01070_),
    .S0(_00357_),
    .S1(net482),
    .X(_01071_));
 sky130_fd_sc_hd__mux4_2 _42000_ (.A0(_01046_),
    .A1(_01047_),
    .A2(_01048_),
    .A3(_01049_),
    .S0(_00357_),
    .S1(net481),
    .X(_01050_));
 sky130_fd_sc_hd__mux4_1 _42001_ (.A0(_01051_),
    .A1(_01052_),
    .A2(_01053_),
    .A3(_01054_),
    .S0(_00357_),
    .S1(net481),
    .X(_01055_));
 sky130_fd_sc_hd__mux4_1 _42002_ (.A0(_01056_),
    .A1(_01057_),
    .A2(_01058_),
    .A3(_01059_),
    .S0(_00357_),
    .S1(net482),
    .X(_01060_));
 sky130_fd_sc_hd__mux4_2 _42003_ (.A0(_01061_),
    .A1(_01062_),
    .A2(_01063_),
    .A3(_01064_),
    .S0(_00357_),
    .S1(net481),
    .X(_01065_));
 sky130_fd_sc_hd__mux4_2 _42004_ (.A0(_01050_),
    .A1(_01055_),
    .A2(_01060_),
    .A3(_01065_),
    .S0(net490),
    .S1(net493),
    .X(_01066_));
 sky130_fd_sc_hd__mux4_2 _42005_ (.A0(_01040_),
    .A1(_01041_),
    .A2(_01042_),
    .A3(_01043_),
    .S0(_00357_),
    .S1(net483),
    .X(_01044_));
 sky130_fd_sc_hd__mux4_2 _42006_ (.A0(_01019_),
    .A1(_01020_),
    .A2(_01021_),
    .A3(_01022_),
    .S0(_00357_),
    .S1(net482),
    .X(_01023_));
 sky130_fd_sc_hd__mux4_2 _42007_ (.A0(_01024_),
    .A1(_01025_),
    .A2(_01026_),
    .A3(_01027_),
    .S0(_00357_),
    .S1(net483),
    .X(_01028_));
 sky130_fd_sc_hd__mux4_1 _42008_ (.A0(_01029_),
    .A1(_01030_),
    .A2(_01031_),
    .A3(_01032_),
    .S0(_00357_),
    .S1(net483),
    .X(_01033_));
 sky130_fd_sc_hd__mux4_2 _42009_ (.A0(_01034_),
    .A1(_01035_),
    .A2(_01036_),
    .A3(_01037_),
    .S0(_00357_),
    .S1(net482),
    .X(_01038_));
 sky130_fd_sc_hd__mux4_1 _42010_ (.A0(_01023_),
    .A1(_01028_),
    .A2(_01033_),
    .A3(_01038_),
    .S0(net490),
    .S1(net493),
    .X(_01039_));
 sky130_fd_sc_hd__mux4_2 _42011_ (.A0(_01013_),
    .A1(_01014_),
    .A2(_01015_),
    .A3(_01016_),
    .S0(_00357_),
    .S1(net483),
    .X(_01017_));
 sky130_fd_sc_hd__mux4_2 _42012_ (.A0(_00992_),
    .A1(_00993_),
    .A2(_00994_),
    .A3(_00995_),
    .S0(_00357_),
    .S1(net482),
    .X(_00996_));
 sky130_fd_sc_hd__mux4_2 _42013_ (.A0(_00997_),
    .A1(_00998_),
    .A2(_00999_),
    .A3(_01000_),
    .S0(_00357_),
    .S1(net483),
    .X(_01001_));
 sky130_fd_sc_hd__mux4_1 _42014_ (.A0(_01002_),
    .A1(_01003_),
    .A2(_01004_),
    .A3(_01005_),
    .S0(_00357_),
    .S1(net483),
    .X(_01006_));
 sky130_fd_sc_hd__mux4_2 _42015_ (.A0(_01007_),
    .A1(_01008_),
    .A2(_01009_),
    .A3(_01010_),
    .S0(_00357_),
    .S1(net482),
    .X(_01011_));
 sky130_fd_sc_hd__mux4_1 _42016_ (.A0(_00996_),
    .A1(_01001_),
    .A2(_01006_),
    .A3(_01011_),
    .S0(net490),
    .S1(net493),
    .X(_01012_));
 sky130_fd_sc_hd__mux4_2 _42017_ (.A0(_00986_),
    .A1(_00987_),
    .A2(_00988_),
    .A3(_00989_),
    .S0(_00357_),
    .S1(net483),
    .X(_00990_));
 sky130_fd_sc_hd__mux4_2 _42018_ (.A0(_00965_),
    .A1(_00966_),
    .A2(_00967_),
    .A3(_00968_),
    .S0(_00357_),
    .S1(net482),
    .X(_00969_));
 sky130_fd_sc_hd__mux4_2 _42019_ (.A0(_00970_),
    .A1(_00971_),
    .A2(_00972_),
    .A3(_00973_),
    .S0(_00357_),
    .S1(net483),
    .X(_00974_));
 sky130_fd_sc_hd__mux4_1 _42020_ (.A0(_00975_),
    .A1(_00976_),
    .A2(_00977_),
    .A3(_00978_),
    .S0(_00357_),
    .S1(net483),
    .X(_00979_));
 sky130_fd_sc_hd__mux4_2 _42021_ (.A0(_00980_),
    .A1(_00981_),
    .A2(_00982_),
    .A3(_00983_),
    .S0(_00357_),
    .S1(net482),
    .X(_00984_));
 sky130_fd_sc_hd__mux4_2 _42022_ (.A0(_00969_),
    .A1(_00974_),
    .A2(_00979_),
    .A3(_00984_),
    .S0(net490),
    .S1(net493),
    .X(_00985_));
 sky130_fd_sc_hd__mux4_2 _42023_ (.A0(_00959_),
    .A1(_00960_),
    .A2(_00961_),
    .A3(_00962_),
    .S0(_00357_),
    .S1(net483),
    .X(_00963_));
 sky130_fd_sc_hd__mux4_2 _42024_ (.A0(_00938_),
    .A1(_00939_),
    .A2(_00940_),
    .A3(_00941_),
    .S0(_00357_),
    .S1(net482),
    .X(_00942_));
 sky130_fd_sc_hd__mux4_2 _42025_ (.A0(_00943_),
    .A1(_00944_),
    .A2(_00945_),
    .A3(_00946_),
    .S0(_00357_),
    .S1(net483),
    .X(_00947_));
 sky130_fd_sc_hd__mux4_1 _42026_ (.A0(_00948_),
    .A1(_00949_),
    .A2(_00950_),
    .A3(_00951_),
    .S0(_00357_),
    .S1(net483),
    .X(_00952_));
 sky130_fd_sc_hd__mux4_1 _42027_ (.A0(_00953_),
    .A1(_00954_),
    .A2(_00955_),
    .A3(_00956_),
    .S0(_00357_),
    .S1(net482),
    .X(_00957_));
 sky130_fd_sc_hd__mux4_1 _42028_ (.A0(_00942_),
    .A1(_00947_),
    .A2(_00952_),
    .A3(_00957_),
    .S0(net490),
    .S1(net493),
    .X(_00958_));
 sky130_fd_sc_hd__mux4_2 _42029_ (.A0(_00932_),
    .A1(_00933_),
    .A2(_00934_),
    .A3(_00935_),
    .S0(_00357_),
    .S1(net483),
    .X(_00936_));
 sky130_fd_sc_hd__mux4_2 _42030_ (.A0(_00911_),
    .A1(_00912_),
    .A2(_00913_),
    .A3(_00914_),
    .S0(_00357_),
    .S1(net482),
    .X(_00915_));
 sky130_fd_sc_hd__mux4_2 _42031_ (.A0(_00916_),
    .A1(_00917_),
    .A2(_00918_),
    .A3(_00919_),
    .S0(_00357_),
    .S1(net483),
    .X(_00920_));
 sky130_fd_sc_hd__mux4_1 _42032_ (.A0(_00921_),
    .A1(_00922_),
    .A2(_00923_),
    .A3(_00924_),
    .S0(_00357_),
    .S1(net483),
    .X(_00925_));
 sky130_fd_sc_hd__mux4_2 _42033_ (.A0(_00926_),
    .A1(_00927_),
    .A2(_00928_),
    .A3(_00929_),
    .S0(_00357_),
    .S1(net482),
    .X(_00930_));
 sky130_fd_sc_hd__mux4_1 _42034_ (.A0(_00915_),
    .A1(_00920_),
    .A2(_00925_),
    .A3(_00930_),
    .S0(net490),
    .S1(net493),
    .X(_00931_));
 sky130_fd_sc_hd__mux4_2 _42035_ (.A0(_00905_),
    .A1(_00906_),
    .A2(_00907_),
    .A3(_00908_),
    .S0(_00357_),
    .S1(net483),
    .X(_00909_));
 sky130_fd_sc_hd__mux4_2 _42036_ (.A0(_00884_),
    .A1(_00885_),
    .A2(_00886_),
    .A3(_00887_),
    .S0(_00357_),
    .S1(net482),
    .X(_00888_));
 sky130_fd_sc_hd__mux4_2 _42037_ (.A0(_00889_),
    .A1(_00890_),
    .A2(_00891_),
    .A3(_00892_),
    .S0(_00357_),
    .S1(net483),
    .X(_00893_));
 sky130_fd_sc_hd__mux4_1 _42038_ (.A0(_00894_),
    .A1(_00895_),
    .A2(_00896_),
    .A3(_00897_),
    .S0(_00357_),
    .S1(net482),
    .X(_00898_));
 sky130_fd_sc_hd__mux4_1 _42039_ (.A0(_00899_),
    .A1(_00900_),
    .A2(_00901_),
    .A3(_00902_),
    .S0(_00357_),
    .S1(net482),
    .X(_00903_));
 sky130_fd_sc_hd__mux4_1 _42040_ (.A0(_00888_),
    .A1(_00893_),
    .A2(_00898_),
    .A3(_00903_),
    .S0(net490),
    .S1(net493),
    .X(_00904_));
 sky130_fd_sc_hd__mux4_2 _42041_ (.A0(_00878_),
    .A1(_00879_),
    .A2(_00880_),
    .A3(_00881_),
    .S0(_00357_),
    .S1(net488),
    .X(_00882_));
 sky130_fd_sc_hd__mux4_2 _42042_ (.A0(_00857_),
    .A1(_00858_),
    .A2(_00859_),
    .A3(_00860_),
    .S0(_00357_),
    .S1(net488),
    .X(_00861_));
 sky130_fd_sc_hd__mux4_2 _42043_ (.A0(_00862_),
    .A1(_00863_),
    .A2(_00864_),
    .A3(_00865_),
    .S0(_00357_),
    .S1(net488),
    .X(_00866_));
 sky130_fd_sc_hd__mux4_2 _42044_ (.A0(_00867_),
    .A1(_00868_),
    .A2(_00869_),
    .A3(_00870_),
    .S0(_00357_),
    .S1(net488),
    .X(_00871_));
 sky130_fd_sc_hd__mux4_1 _42045_ (.A0(_00872_),
    .A1(_00873_),
    .A2(_00874_),
    .A3(_00875_),
    .S0(_00357_),
    .S1(net488),
    .X(_00876_));
 sky130_fd_sc_hd__mux4_2 _42046_ (.A0(_00861_),
    .A1(_00866_),
    .A2(_00871_),
    .A3(_00876_),
    .S0(net491),
    .S1(net493),
    .X(_00877_));
 sky130_fd_sc_hd__mux4_2 _42047_ (.A0(_00851_),
    .A1(_00852_),
    .A2(_00853_),
    .A3(_00854_),
    .S0(_00357_),
    .S1(net488),
    .X(_00855_));
 sky130_fd_sc_hd__mux4_2 _42048_ (.A0(_00830_),
    .A1(_00831_),
    .A2(_00832_),
    .A3(_00833_),
    .S0(net480),
    .S1(net487),
    .X(_00834_));
 sky130_fd_sc_hd__mux4_2 _42049_ (.A0(_00835_),
    .A1(_00836_),
    .A2(_00837_),
    .A3(_00838_),
    .S0(_00357_),
    .S1(net488),
    .X(_00839_));
 sky130_fd_sc_hd__mux4_2 _42050_ (.A0(_00840_),
    .A1(_00841_),
    .A2(_00842_),
    .A3(_00843_),
    .S0(net480),
    .S1(net487),
    .X(_00844_));
 sky130_fd_sc_hd__mux4_1 _42051_ (.A0(_00845_),
    .A1(_00846_),
    .A2(_00847_),
    .A3(_00848_),
    .S0(net480),
    .S1(net487),
    .X(_00849_));
 sky130_fd_sc_hd__mux4_2 _42052_ (.A0(_00834_),
    .A1(_00839_),
    .A2(_00844_),
    .A3(_00849_),
    .S0(net491),
    .S1(net492),
    .X(_00850_));
 sky130_fd_sc_hd__mux4_1 _42053_ (.A0(_00824_),
    .A1(_00825_),
    .A2(_00826_),
    .A3(_00827_),
    .S0(net480),
    .S1(net487),
    .X(_00828_));
 sky130_fd_sc_hd__mux4_2 _42054_ (.A0(_00803_),
    .A1(_00804_),
    .A2(_00805_),
    .A3(_00806_),
    .S0(net480),
    .S1(net487),
    .X(_00807_));
 sky130_fd_sc_hd__mux4_1 _42055_ (.A0(_00808_),
    .A1(_00809_),
    .A2(_00810_),
    .A3(_00811_),
    .S0(net480),
    .S1(net487),
    .X(_00812_));
 sky130_fd_sc_hd__mux4_2 _42056_ (.A0(_00813_),
    .A1(_00814_),
    .A2(_00815_),
    .A3(_00816_),
    .S0(net480),
    .S1(net487),
    .X(_00817_));
 sky130_fd_sc_hd__mux4_1 _42057_ (.A0(_00818_),
    .A1(_00819_),
    .A2(_00820_),
    .A3(_00821_),
    .S0(net480),
    .S1(net487),
    .X(_00822_));
 sky130_fd_sc_hd__mux4_2 _42058_ (.A0(_00807_),
    .A1(_00812_),
    .A2(_00817_),
    .A3(_00822_),
    .S0(net491),
    .S1(net492),
    .X(_00823_));
 sky130_fd_sc_hd__mux4_2 _42059_ (.A0(_00797_),
    .A1(_00798_),
    .A2(_00799_),
    .A3(_00800_),
    .S0(net480),
    .S1(net488),
    .X(_00801_));
 sky130_fd_sc_hd__mux4_2 _42060_ (.A0(_00776_),
    .A1(_00777_),
    .A2(_00778_),
    .A3(_00779_),
    .S0(net480),
    .S1(net487),
    .X(_00780_));
 sky130_fd_sc_hd__mux4_2 _42061_ (.A0(_00781_),
    .A1(_00782_),
    .A2(_00783_),
    .A3(_00784_),
    .S0(net480),
    .S1(net488),
    .X(_00785_));
 sky130_fd_sc_hd__mux4_1 _42062_ (.A0(_00786_),
    .A1(_00787_),
    .A2(_00788_),
    .A3(_00789_),
    .S0(net480),
    .S1(net487),
    .X(_00790_));
 sky130_fd_sc_hd__mux4_1 _42063_ (.A0(_00791_),
    .A1(_00792_),
    .A2(_00793_),
    .A3(_00794_),
    .S0(net480),
    .S1(net487),
    .X(_00795_));
 sky130_fd_sc_hd__mux4_2 _42064_ (.A0(_00780_),
    .A1(_00785_),
    .A2(_00790_),
    .A3(_00795_),
    .S0(net491),
    .S1(net492),
    .X(_00796_));
 sky130_fd_sc_hd__mux4_1 _42065_ (.A0(_00770_),
    .A1(_00771_),
    .A2(_00772_),
    .A3(_00773_),
    .S0(net480),
    .S1(net487),
    .X(_00774_));
 sky130_fd_sc_hd__mux4_2 _42066_ (.A0(_00749_),
    .A1(_00750_),
    .A2(_00751_),
    .A3(_00752_),
    .S0(net480),
    .S1(net487),
    .X(_00753_));
 sky130_fd_sc_hd__mux4_1 _42067_ (.A0(_00754_),
    .A1(_00755_),
    .A2(_00756_),
    .A3(_00757_),
    .S0(net480),
    .S1(net487),
    .X(_00758_));
 sky130_fd_sc_hd__mux4_1 _42068_ (.A0(_00759_),
    .A1(_00760_),
    .A2(_00761_),
    .A3(_00762_),
    .S0(net480),
    .S1(net487),
    .X(_00763_));
 sky130_fd_sc_hd__mux4_1 _42069_ (.A0(_00764_),
    .A1(_00765_),
    .A2(_00766_),
    .A3(_00767_),
    .S0(net480),
    .S1(net487),
    .X(_00768_));
 sky130_fd_sc_hd__mux4_2 _42070_ (.A0(_00753_),
    .A1(_00758_),
    .A2(_00763_),
    .A3(_00768_),
    .S0(net491),
    .S1(net492),
    .X(_00769_));
 sky130_fd_sc_hd__mux4_1 _42071_ (.A0(_00743_),
    .A1(_00744_),
    .A2(_00745_),
    .A3(_00746_),
    .S0(net480),
    .S1(net487),
    .X(_00747_));
 sky130_fd_sc_hd__mux4_1 _42072_ (.A0(_00722_),
    .A1(_00723_),
    .A2(_00724_),
    .A3(_00725_),
    .S0(net480),
    .S1(net486),
    .X(_00726_));
 sky130_fd_sc_hd__mux4_2 _42073_ (.A0(_00727_),
    .A1(_00728_),
    .A2(_00729_),
    .A3(_00730_),
    .S0(net480),
    .S1(net486),
    .X(_00731_));
 sky130_fd_sc_hd__mux4_1 _42074_ (.A0(_00732_),
    .A1(_00733_),
    .A2(_00734_),
    .A3(_00735_),
    .S0(net480),
    .S1(net486),
    .X(_00736_));
 sky130_fd_sc_hd__mux4_2 _42075_ (.A0(_00737_),
    .A1(_00738_),
    .A2(_00739_),
    .A3(_00740_),
    .S0(net480),
    .S1(net487),
    .X(_00741_));
 sky130_fd_sc_hd__mux4_2 _42076_ (.A0(_00726_),
    .A1(_00731_),
    .A2(_00736_),
    .A3(_00741_),
    .S0(net491),
    .S1(net492),
    .X(_00742_));
 sky130_fd_sc_hd__mux4_1 _42077_ (.A0(_00716_),
    .A1(_00717_),
    .A2(_00718_),
    .A3(_00719_),
    .S0(net480),
    .S1(net486),
    .X(_00720_));
 sky130_fd_sc_hd__mux4_2 _42078_ (.A0(_00695_),
    .A1(_00696_),
    .A2(_00697_),
    .A3(_00698_),
    .S0(net480),
    .S1(net486),
    .X(_00699_));
 sky130_fd_sc_hd__mux4_2 _42079_ (.A0(_00700_),
    .A1(_00701_),
    .A2(_00702_),
    .A3(_00703_),
    .S0(net480),
    .S1(net486),
    .X(_00704_));
 sky130_fd_sc_hd__mux4_1 _42080_ (.A0(_00705_),
    .A1(_00706_),
    .A2(_00707_),
    .A3(_00708_),
    .S0(net480),
    .S1(net486),
    .X(_00709_));
 sky130_fd_sc_hd__mux4_2 _42081_ (.A0(_00710_),
    .A1(_00711_),
    .A2(_00712_),
    .A3(_00713_),
    .S0(net480),
    .S1(net486),
    .X(_00714_));
 sky130_fd_sc_hd__mux4_2 _42082_ (.A0(_00699_),
    .A1(_00704_),
    .A2(_00709_),
    .A3(_00714_),
    .S0(net489),
    .S1(net492),
    .X(_00715_));
 sky130_fd_sc_hd__mux4_1 _42083_ (.A0(_00689_),
    .A1(_00690_),
    .A2(_00691_),
    .A3(_00692_),
    .S0(net480),
    .S1(net486),
    .X(_00693_));
 sky130_fd_sc_hd__mux4_2 _42084_ (.A0(_00668_),
    .A1(_00669_),
    .A2(_00670_),
    .A3(_00671_),
    .S0(net480),
    .S1(net486),
    .X(_00672_));
 sky130_fd_sc_hd__mux4_2 _42085_ (.A0(_00673_),
    .A1(_00674_),
    .A2(_00675_),
    .A3(_00676_),
    .S0(net480),
    .S1(net486),
    .X(_00677_));
 sky130_fd_sc_hd__mux4_1 _42086_ (.A0(_00678_),
    .A1(_00679_),
    .A2(_00680_),
    .A3(_00681_),
    .S0(net480),
    .S1(net486),
    .X(_00682_));
 sky130_fd_sc_hd__mux4_1 _42087_ (.A0(_00683_),
    .A1(_00684_),
    .A2(_00685_),
    .A3(_00686_),
    .S0(net480),
    .S1(net486),
    .X(_00687_));
 sky130_fd_sc_hd__mux4_2 _42088_ (.A0(_00672_),
    .A1(_00677_),
    .A2(_00682_),
    .A3(_00687_),
    .S0(net489),
    .S1(net492),
    .X(_00688_));
 sky130_fd_sc_hd__mux4_2 _42089_ (.A0(_00662_),
    .A1(_00663_),
    .A2(_00664_),
    .A3(_00665_),
    .S0(net480),
    .S1(net485),
    .X(_00666_));
 sky130_fd_sc_hd__mux4_2 _42090_ (.A0(_00641_),
    .A1(_00642_),
    .A2(_00643_),
    .A3(_00644_),
    .S0(net480),
    .S1(net485),
    .X(_00645_));
 sky130_fd_sc_hd__mux4_2 _42091_ (.A0(_00646_),
    .A1(_00647_),
    .A2(_00648_),
    .A3(_00649_),
    .S0(net480),
    .S1(net485),
    .X(_00650_));
 sky130_fd_sc_hd__mux4_1 _42092_ (.A0(_00651_),
    .A1(_00652_),
    .A2(_00653_),
    .A3(_00654_),
    .S0(net480),
    .S1(net485),
    .X(_00655_));
 sky130_fd_sc_hd__mux4_1 _42093_ (.A0(_00656_),
    .A1(_00657_),
    .A2(_00658_),
    .A3(_00659_),
    .S0(net480),
    .S1(net485),
    .X(_00660_));
 sky130_fd_sc_hd__mux4_2 _42094_ (.A0(_00645_),
    .A1(_00650_),
    .A2(_00655_),
    .A3(_00660_),
    .S0(net489),
    .S1(net492),
    .X(_00661_));
 sky130_fd_sc_hd__mux4_2 _42095_ (.A0(_00635_),
    .A1(_00636_),
    .A2(_00637_),
    .A3(_00638_),
    .S0(net480),
    .S1(net485),
    .X(_00639_));
 sky130_fd_sc_hd__mux4_2 _42096_ (.A0(_00614_),
    .A1(_00615_),
    .A2(_00616_),
    .A3(_00617_),
    .S0(net480),
    .S1(net485),
    .X(_00618_));
 sky130_fd_sc_hd__mux4_2 _42097_ (.A0(_00619_),
    .A1(_00620_),
    .A2(_00621_),
    .A3(_00622_),
    .S0(net480),
    .S1(net485),
    .X(_00623_));
 sky130_fd_sc_hd__mux4_1 _42098_ (.A0(_00624_),
    .A1(_00625_),
    .A2(_00626_),
    .A3(_00627_),
    .S0(net480),
    .S1(net485),
    .X(_00628_));
 sky130_fd_sc_hd__mux4_2 _42099_ (.A0(_00629_),
    .A1(_00630_),
    .A2(_00631_),
    .A3(_00632_),
    .S0(net480),
    .S1(net485),
    .X(_00633_));
 sky130_fd_sc_hd__mux4_2 _42100_ (.A0(_00618_),
    .A1(_00623_),
    .A2(_00628_),
    .A3(_00633_),
    .S0(net489),
    .S1(net492),
    .X(_00634_));
 sky130_fd_sc_hd__mux4_1 _42101_ (.A0(_00608_),
    .A1(_00609_),
    .A2(_00610_),
    .A3(_00611_),
    .S0(net480),
    .S1(net486),
    .X(_00612_));
 sky130_fd_sc_hd__mux4_2 _42102_ (.A0(_00587_),
    .A1(_00588_),
    .A2(_00589_),
    .A3(_00590_),
    .S0(net480),
    .S1(net486),
    .X(_00591_));
 sky130_fd_sc_hd__mux4_2 _42103_ (.A0(_00592_),
    .A1(_00593_),
    .A2(_00594_),
    .A3(_00595_),
    .S0(net480),
    .S1(net486),
    .X(_00596_));
 sky130_fd_sc_hd__mux4_1 _42104_ (.A0(_00597_),
    .A1(_00598_),
    .A2(_00599_),
    .A3(_00600_),
    .S0(net480),
    .S1(net486),
    .X(_00601_));
 sky130_fd_sc_hd__mux4_2 _42105_ (.A0(_00602_),
    .A1(_00603_),
    .A2(_00604_),
    .A3(_00605_),
    .S0(net480),
    .S1(net486),
    .X(_00606_));
 sky130_fd_sc_hd__mux4_2 _42106_ (.A0(_00591_),
    .A1(_00596_),
    .A2(_00601_),
    .A3(_00606_),
    .S0(net489),
    .S1(net492),
    .X(_00607_));
 sky130_fd_sc_hd__mux4_1 _42107_ (.A0(_00581_),
    .A1(_00582_),
    .A2(_00583_),
    .A3(_00584_),
    .S0(net480),
    .S1(net486),
    .X(_00585_));
 sky130_fd_sc_hd__mux4_2 _42108_ (.A0(_00560_),
    .A1(_00561_),
    .A2(_00562_),
    .A3(_00563_),
    .S0(net480),
    .S1(net486),
    .X(_00564_));
 sky130_fd_sc_hd__mux4_2 _42109_ (.A0(_00565_),
    .A1(_00566_),
    .A2(_00567_),
    .A3(_00568_),
    .S0(net480),
    .S1(net486),
    .X(_00569_));
 sky130_fd_sc_hd__mux4_1 _42110_ (.A0(_00570_),
    .A1(_00571_),
    .A2(_00572_),
    .A3(_00573_),
    .S0(net480),
    .S1(net485),
    .X(_00574_));
 sky130_fd_sc_hd__mux4_1 _42111_ (.A0(_00575_),
    .A1(_00576_),
    .A2(_00577_),
    .A3(_00578_),
    .S0(net480),
    .S1(net485),
    .X(_00579_));
 sky130_fd_sc_hd__mux4_2 _42112_ (.A0(_00564_),
    .A1(_00569_),
    .A2(_00574_),
    .A3(_00579_),
    .S0(net489),
    .S1(net492),
    .X(_00580_));
 sky130_fd_sc_hd__mux4_1 _42113_ (.A0(_00554_),
    .A1(_00555_),
    .A2(_00556_),
    .A3(_00557_),
    .S0(net480),
    .S1(net484),
    .X(_00558_));
 sky130_fd_sc_hd__mux4_2 _42114_ (.A0(_00533_),
    .A1(_00534_),
    .A2(_00535_),
    .A3(_00536_),
    .S0(net480),
    .S1(net485),
    .X(_00537_));
 sky130_fd_sc_hd__mux4_1 _42115_ (.A0(_00538_),
    .A1(_00539_),
    .A2(_00540_),
    .A3(_00541_),
    .S0(net480),
    .S1(net485),
    .X(_00542_));
 sky130_fd_sc_hd__mux4_2 _42116_ (.A0(_00543_),
    .A1(_00544_),
    .A2(_00545_),
    .A3(_00546_),
    .S0(net480),
    .S1(net485),
    .X(_00547_));
 sky130_fd_sc_hd__mux4_1 _42117_ (.A0(_00548_),
    .A1(_00549_),
    .A2(_00550_),
    .A3(_00551_),
    .S0(net480),
    .S1(net485),
    .X(_00552_));
 sky130_fd_sc_hd__mux4_2 _42118_ (.A0(_00537_),
    .A1(_00542_),
    .A2(_00547_),
    .A3(_00552_),
    .S0(net489),
    .S1(net492),
    .X(_00553_));
 sky130_fd_sc_hd__mux4_2 _42119_ (.A0(_00527_),
    .A1(_00528_),
    .A2(_00529_),
    .A3(_00530_),
    .S0(net480),
    .S1(net484),
    .X(_00531_));
 sky130_fd_sc_hd__mux4_2 _42120_ (.A0(_00506_),
    .A1(_00507_),
    .A2(_00508_),
    .A3(_00509_),
    .S0(net480),
    .S1(net485),
    .X(_00510_));
 sky130_fd_sc_hd__mux4_2 _42121_ (.A0(_00511_),
    .A1(_00512_),
    .A2(_00513_),
    .A3(_00514_),
    .S0(net480),
    .S1(net484),
    .X(_00515_));
 sky130_fd_sc_hd__mux4_1 _42122_ (.A0(_00516_),
    .A1(_00517_),
    .A2(_00518_),
    .A3(_00519_),
    .S0(net480),
    .S1(net484),
    .X(_00520_));
 sky130_fd_sc_hd__mux4_1 _42123_ (.A0(_00521_),
    .A1(_00522_),
    .A2(_00523_),
    .A3(_00524_),
    .S0(net480),
    .S1(net484),
    .X(_00525_));
 sky130_fd_sc_hd__mux4_2 _42124_ (.A0(_00510_),
    .A1(_00515_),
    .A2(_00520_),
    .A3(_00525_),
    .S0(net489),
    .S1(net492),
    .X(_00526_));
 sky130_fd_sc_hd__mux4_1 _42125_ (.A0(_00500_),
    .A1(_00501_),
    .A2(_00502_),
    .A3(_00503_),
    .S0(net480),
    .S1(net484),
    .X(_00504_));
 sky130_fd_sc_hd__mux4_2 _42126_ (.A0(_00479_),
    .A1(_00480_),
    .A2(_00481_),
    .A3(_00482_),
    .S0(net480),
    .S1(net485),
    .X(_00483_));
 sky130_fd_sc_hd__mux4_1 _42127_ (.A0(_00484_),
    .A1(_00485_),
    .A2(_00486_),
    .A3(_00487_),
    .S0(net480),
    .S1(net484),
    .X(_00488_));
 sky130_fd_sc_hd__mux4_2 _42128_ (.A0(_00489_),
    .A1(_00490_),
    .A2(_00491_),
    .A3(_00492_),
    .S0(net480),
    .S1(net485),
    .X(_00493_));
 sky130_fd_sc_hd__mux4_1 _42129_ (.A0(_00494_),
    .A1(_00495_),
    .A2(_00496_),
    .A3(_00497_),
    .S0(net480),
    .S1(net485),
    .X(_00498_));
 sky130_fd_sc_hd__mux4_2 _42130_ (.A0(_00483_),
    .A1(_00488_),
    .A2(_00493_),
    .A3(_00498_),
    .S0(net489),
    .S1(net492),
    .X(_00499_));
 sky130_fd_sc_hd__mux4_2 _42131_ (.A0(_00473_),
    .A1(_00474_),
    .A2(_00475_),
    .A3(_00476_),
    .S0(net480),
    .S1(net484),
    .X(_00477_));
 sky130_fd_sc_hd__mux4_1 _42132_ (.A0(_00452_),
    .A1(_00453_),
    .A2(_00454_),
    .A3(_00455_),
    .S0(net480),
    .S1(net484),
    .X(_00456_));
 sky130_fd_sc_hd__mux4_2 _42133_ (.A0(_00457_),
    .A1(_00458_),
    .A2(_00459_),
    .A3(_00460_),
    .S0(net480),
    .S1(net484),
    .X(_00461_));
 sky130_fd_sc_hd__mux4_1 _42134_ (.A0(_00462_),
    .A1(_00463_),
    .A2(_00464_),
    .A3(_00465_),
    .S0(net480),
    .S1(net484),
    .X(_00466_));
 sky130_fd_sc_hd__mux4_2 _42135_ (.A0(_00467_),
    .A1(_00468_),
    .A2(_00469_),
    .A3(_00470_),
    .S0(net480),
    .S1(net484),
    .X(_00471_));
 sky130_fd_sc_hd__mux4_2 _42136_ (.A0(_00456_),
    .A1(_00461_),
    .A2(_00466_),
    .A3(_00471_),
    .S0(net489),
    .S1(net492),
    .X(_00472_));
 sky130_fd_sc_hd__mux4_2 _42137_ (.A0(_00446_),
    .A1(_00447_),
    .A2(_00448_),
    .A3(_00449_),
    .S0(net480),
    .S1(net484),
    .X(_00450_));
 sky130_fd_sc_hd__mux4_1 _42138_ (.A0(_00425_),
    .A1(_00426_),
    .A2(_00427_),
    .A3(_00428_),
    .S0(net480),
    .S1(net484),
    .X(_00429_));
 sky130_fd_sc_hd__mux4_1 _42139_ (.A0(_00430_),
    .A1(_00431_),
    .A2(_00432_),
    .A3(_00433_),
    .S0(net480),
    .S1(net484),
    .X(_00434_));
 sky130_fd_sc_hd__mux4_1 _42140_ (.A0(_00435_),
    .A1(_00436_),
    .A2(_00437_),
    .A3(_00438_),
    .S0(net480),
    .S1(net484),
    .X(_00439_));
 sky130_fd_sc_hd__mux4_2 _42141_ (.A0(_00440_),
    .A1(_00441_),
    .A2(_00442_),
    .A3(_00443_),
    .S0(net480),
    .S1(net484),
    .X(_00444_));
 sky130_fd_sc_hd__mux4_2 _42142_ (.A0(_00429_),
    .A1(_00434_),
    .A2(_00439_),
    .A3(_00444_),
    .S0(net489),
    .S1(net492),
    .X(_00445_));
 sky130_fd_sc_hd__mux4_1 _42143_ (.A0(_00419_),
    .A1(_00420_),
    .A2(_00421_),
    .A3(_00422_),
    .S0(net480),
    .S1(net484),
    .X(_00423_));
 sky130_fd_sc_hd__mux4_2 _42144_ (.A0(_00398_),
    .A1(_00399_),
    .A2(_00400_),
    .A3(_00401_),
    .S0(net480),
    .S1(net484),
    .X(_00402_));
 sky130_fd_sc_hd__mux4_1 _42145_ (.A0(_00403_),
    .A1(_00404_),
    .A2(_00405_),
    .A3(_00406_),
    .S0(net480),
    .S1(net484),
    .X(_00407_));
 sky130_fd_sc_hd__mux4_2 _42146_ (.A0(_00408_),
    .A1(_00409_),
    .A2(_00410_),
    .A3(_00411_),
    .S0(net480),
    .S1(net484),
    .X(_00412_));
 sky130_fd_sc_hd__mux4_1 _42147_ (.A0(_00413_),
    .A1(_00414_),
    .A2(_00415_),
    .A3(_00416_),
    .S0(net480),
    .S1(net484),
    .X(_00417_));
 sky130_fd_sc_hd__mux4_2 _42148_ (.A0(_00402_),
    .A1(_00407_),
    .A2(_00412_),
    .A3(_00417_),
    .S0(net489),
    .S1(net492),
    .X(_00418_));
 sky130_fd_sc_hd__mux4_1 _42149_ (.A0(_00392_),
    .A1(_00393_),
    .A2(_00394_),
    .A3(_00395_),
    .S0(_00357_),
    .S1(net488),
    .X(_00396_));
 sky130_fd_sc_hd__mux4_2 _42150_ (.A0(_00371_),
    .A1(_00372_),
    .A2(_00373_),
    .A3(_00374_),
    .S0(_00357_),
    .S1(net488),
    .X(_00375_));
 sky130_fd_sc_hd__mux4_2 _42151_ (.A0(_00376_),
    .A1(_00377_),
    .A2(_00378_),
    .A3(_00379_),
    .S0(_00357_),
    .S1(net488),
    .X(_00380_));
 sky130_fd_sc_hd__mux4_1 _42152_ (.A0(_00381_),
    .A1(_00382_),
    .A2(_00383_),
    .A3(_00384_),
    .S0(_00357_),
    .S1(net488),
    .X(_00385_));
 sky130_fd_sc_hd__mux4_1 _42153_ (.A0(_00386_),
    .A1(_00387_),
    .A2(_00388_),
    .A3(_00389_),
    .S0(_00357_),
    .S1(net488),
    .X(_00390_));
 sky130_fd_sc_hd__mux4_2 _42154_ (.A0(_00375_),
    .A1(_00380_),
    .A2(_00385_),
    .A3(_00390_),
    .S0(net491),
    .S1(net493),
    .X(_00391_));
 sky130_fd_sc_hd__mux4_1 _42155_ (.A0(\cpuregs[16][0] ),
    .A1(\cpuregs[17][0] ),
    .A2(\cpuregs[18][0] ),
    .A3(\cpuregs[19][0] ),
    .S0(_00357_),
    .S1(net483),
    .X(_00369_));
 sky130_fd_sc_hd__mux4_2 _42156_ (.A0(\cpuregs[0][0] ),
    .A1(\cpuregs[1][0] ),
    .A2(\cpuregs[2][0] ),
    .A3(\cpuregs[3][0] ),
    .S0(_00357_),
    .S1(net488),
    .X(_00359_));
 sky130_fd_sc_hd__mux4_2 _42157_ (.A0(\cpuregs[4][0] ),
    .A1(\cpuregs[5][0] ),
    .A2(\cpuregs[6][0] ),
    .A3(\cpuregs[7][0] ),
    .S0(_00357_),
    .S1(net483),
    .X(_00361_));
 sky130_fd_sc_hd__mux4_1 _42158_ (.A0(\cpuregs[8][0] ),
    .A1(\cpuregs[9][0] ),
    .A2(\cpuregs[10][0] ),
    .A3(\cpuregs[11][0] ),
    .S0(_00357_),
    .S1(net488),
    .X(_00363_));
 sky130_fd_sc_hd__mux4_1 _42159_ (.A0(\cpuregs[12][0] ),
    .A1(\cpuregs[13][0] ),
    .A2(\cpuregs[14][0] ),
    .A3(\cpuregs[15][0] ),
    .S0(_00357_),
    .S1(net483),
    .X(_00364_));
 sky130_fd_sc_hd__mux4_2 _42160_ (.A0(_00359_),
    .A1(_00361_),
    .A2(_00363_),
    .A3(_00364_),
    .S0(net490),
    .S1(net493),
    .X(_00365_));
 sky130_fd_sc_hd__mux4_1 _42161_ (.A0(_02581_),
    .A1(_01681_),
    .A2(_01679_),
    .A3(_02581_),
    .S0(net428),
    .S1(_00309_),
    .X(_01682_));
 sky130_fd_sc_hd__mux4_1 _42162_ (.A0(_02580_),
    .A1(_01677_),
    .A2(_01675_),
    .A3(_02580_),
    .S0(net428),
    .S1(_00309_),
    .X(_01678_));
 sky130_fd_sc_hd__mux4_1 _42163_ (.A0(_02579_),
    .A1(_01673_),
    .A2(_01671_),
    .A3(_02579_),
    .S0(net428),
    .S1(_00309_),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_1 _42164_ (.A0(_02578_),
    .A1(_01669_),
    .A2(_01667_),
    .A3(_02578_),
    .S0(net428),
    .S1(_00309_),
    .X(_01670_));
 sky130_fd_sc_hd__mux4_1 _42165_ (.A0(_02577_),
    .A1(_01665_),
    .A2(_01663_),
    .A3(_02577_),
    .S0(net428),
    .S1(_00309_),
    .X(_01666_));
 sky130_fd_sc_hd__mux4_1 _42166_ (.A0(_02576_),
    .A1(_01661_),
    .A2(_01659_),
    .A3(_02576_),
    .S0(net428),
    .S1(_00309_),
    .X(_01662_));
 sky130_fd_sc_hd__mux4_1 _42167_ (.A0(_02575_),
    .A1(_01657_),
    .A2(_01655_),
    .A3(_02575_),
    .S0(net428),
    .S1(_00309_),
    .X(_01658_));
 sky130_fd_sc_hd__mux4_1 _42168_ (.A0(_02574_),
    .A1(_01653_),
    .A2(_01651_),
    .A3(_02574_),
    .S0(net428),
    .S1(_00309_),
    .X(_01654_));
 sky130_fd_sc_hd__mux4_1 _42169_ (.A0(_02573_),
    .A1(_01649_),
    .A2(_01647_),
    .A3(_02573_),
    .S0(net428),
    .S1(_00309_),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_1 _42170_ (.A0(_02572_),
    .A1(_01645_),
    .A2(_01643_),
    .A3(_02572_),
    .S0(net428),
    .S1(_00309_),
    .X(_01646_));
 sky130_fd_sc_hd__mux4_1 _42171_ (.A0(_02570_),
    .A1(_01641_),
    .A2(_01639_),
    .A3(_02570_),
    .S0(net428),
    .S1(_00309_),
    .X(_01642_));
 sky130_fd_sc_hd__mux4_1 _42172_ (.A0(_02569_),
    .A1(_01637_),
    .A2(_01635_),
    .A3(_02569_),
    .S0(net428),
    .S1(_00309_),
    .X(_01638_));
 sky130_fd_sc_hd__mux4_1 _42173_ (.A0(_02568_),
    .A1(_01633_),
    .A2(_01631_),
    .A3(_02568_),
    .S0(net428),
    .S1(_00309_),
    .X(_01634_));
 sky130_fd_sc_hd__mux4_1 _42174_ (.A0(_02567_),
    .A1(_01629_),
    .A2(_01627_),
    .A3(_02567_),
    .S0(net428),
    .S1(_00309_),
    .X(_01630_));
 sky130_fd_sc_hd__mux4_1 _42175_ (.A0(_02566_),
    .A1(_01625_),
    .A2(_01623_),
    .A3(_02566_),
    .S0(net428),
    .S1(_00309_),
    .X(_01626_));
 sky130_fd_sc_hd__mux4_1 _42176_ (.A0(_02565_),
    .A1(_01621_),
    .A2(_01619_),
    .A3(_02565_),
    .S0(net428),
    .S1(_00309_),
    .X(_01622_));
 sky130_fd_sc_hd__mux4_1 _42177_ (.A0(_02564_),
    .A1(_01617_),
    .A2(_01615_),
    .A3(_02564_),
    .S0(net428),
    .S1(_00309_),
    .X(_01618_));
 sky130_fd_sc_hd__mux4_2 _42178_ (.A0(_02563_),
    .A1(_01613_),
    .A2(_01611_),
    .A3(_02563_),
    .S0(net428),
    .S1(_00309_),
    .X(_01614_));
 sky130_fd_sc_hd__mux4_1 _42179_ (.A0(_02562_),
    .A1(_01609_),
    .A2(_01607_),
    .A3(_02562_),
    .S0(net428),
    .S1(_00309_),
    .X(_01610_));
 sky130_fd_sc_hd__mux4_1 _42180_ (.A0(_02561_),
    .A1(_01605_),
    .A2(_01603_),
    .A3(_02561_),
    .S0(net428),
    .S1(_00309_),
    .X(_01606_));
 sky130_fd_sc_hd__mux4_1 _42181_ (.A0(_02589_),
    .A1(_01601_),
    .A2(_01599_),
    .A3(_02589_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01602_));
 sky130_fd_sc_hd__mux4_1 _42182_ (.A0(_02588_),
    .A1(_01597_),
    .A2(_01595_),
    .A3(_02588_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01598_));
 sky130_fd_sc_hd__mux4_1 _42183_ (.A0(_02587_),
    .A1(_01593_),
    .A2(_01591_),
    .A3(_02587_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01594_));
 sky130_fd_sc_hd__mux4_1 _42184_ (.A0(_02586_),
    .A1(_01589_),
    .A2(_01587_),
    .A3(_02586_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _42185_ (.A0(_02585_),
    .A1(_01585_),
    .A2(_01583_),
    .A3(_02585_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01586_));
 sky130_fd_sc_hd__mux4_1 _42186_ (.A0(_02584_),
    .A1(_01581_),
    .A2(_01579_),
    .A3(_02584_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01582_));
 sky130_fd_sc_hd__mux4_1 _42187_ (.A0(_02583_),
    .A1(_01577_),
    .A2(_01575_),
    .A3(_02583_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01578_));
 sky130_fd_sc_hd__mux4_1 _42188_ (.A0(_02582_),
    .A1(_01573_),
    .A2(_01571_),
    .A3(_02582_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01574_));
 sky130_fd_sc_hd__mux4_1 _42189_ (.A0(_02571_),
    .A1(_01569_),
    .A2(_01567_),
    .A3(_02571_),
    .S0(_20894_),
    .S1(_00309_),
    .X(_01570_));
 sky130_fd_sc_hd__dfxtp_1 _42190_ (.D(_02687_),
    .Q(\alu_shl[0] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42191_ (.D(_02688_),
    .Q(\alu_shl[1] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42192_ (.D(_02689_),
    .Q(\alu_shl[2] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42193_ (.D(_02690_),
    .Q(\alu_shl[3] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42194_ (.D(_02691_),
    .Q(\alu_shl[4] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42195_ (.D(_02692_),
    .Q(\alu_shl[5] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42196_ (.D(_02693_),
    .Q(\alu_shl[6] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42197_ (.D(_02694_),
    .Q(\alu_shl[7] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42198_ (.D(_02695_),
    .Q(\alu_shl[8] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42199_ (.D(_02696_),
    .Q(\alu_shl[9] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _42200_ (.D(_02697_),
    .Q(\alu_shl[10] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42201_ (.D(_02698_),
    .Q(\alu_shl[11] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42202_ (.D(_02699_),
    .Q(\alu_shl[12] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42203_ (.D(_02700_),
    .Q(\alu_shl[13] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _42204_ (.D(_02701_),
    .Q(\alu_shl[14] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 _42205_ (.D(_02702_),
    .Q(\alu_shl[15] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_2 _42206_ (.D(_02703_),
    .Q(alu_wait),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _42207_ (.D(_02704_),
    .Q(\latched_rd[3] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 _42208_ (.D(_02705_),
    .Q(\latched_rd[2] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 _42209_ (.D(_02706_),
    .Q(\latched_rd[1] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42210_ (.D(_02707_),
    .Q(\latched_rd[0] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_2 _42211_ (.D(_02708_),
    .Q(\decoded_imm[31] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 _42212_ (.D(_02709_),
    .Q(\decoded_imm[30] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_4 _42213_ (.D(_02710_),
    .Q(\decoded_imm[29] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_2 _42214_ (.D(_02711_),
    .Q(\decoded_imm[28] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _42215_ (.D(_02712_),
    .Q(\decoded_imm[27] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _42216_ (.D(_02713_),
    .Q(\decoded_imm[26] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_2 _42217_ (.D(_02714_),
    .Q(\decoded_imm[25] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 _42218_ (.D(_02715_),
    .Q(\decoded_imm[24] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 _42219_ (.D(_02716_),
    .Q(\decoded_imm[23] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_2 _42220_ (.D(_02717_),
    .Q(\decoded_imm[22] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 _42221_ (.D(_02718_),
    .Q(\decoded_imm[21] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_2 _42222_ (.D(_02719_),
    .Q(\decoded_imm[20] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_2 _42223_ (.D(_02720_),
    .Q(\decoded_imm[19] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42224_ (.D(_02721_),
    .Q(\decoded_imm[18] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42225_ (.D(_02722_),
    .Q(\decoded_imm[17] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 _42226_ (.D(_02723_),
    .Q(\decoded_imm[16] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_2 _42227_ (.D(_02724_),
    .Q(\decoded_imm[15] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_1 _42228_ (.D(_02725_),
    .Q(\decoded_imm[14] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_2 _42229_ (.D(_02726_),
    .Q(\decoded_imm[13] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 _42230_ (.D(_02727_),
    .Q(\decoded_imm[12] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_2 _42231_ (.D(_02728_),
    .Q(\decoded_imm[11] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_2 _42232_ (.D(_02729_),
    .Q(\decoded_imm[10] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42233_ (.D(_02730_),
    .Q(\decoded_imm[9] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _42234_ (.D(_02731_),
    .Q(\decoded_imm[8] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42235_ (.D(_02732_),
    .Q(\decoded_imm[7] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42236_ (.D(_02733_),
    .Q(\decoded_imm[6] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_2 _42237_ (.D(_02734_),
    .Q(\decoded_imm[5] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42238_ (.D(_02735_),
    .Q(\decoded_imm[4] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 _42239_ (.D(_02736_),
    .Q(\decoded_imm[3] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_2 _42240_ (.D(_02737_),
    .Q(\decoded_imm[2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_2 _42241_ (.D(_02738_),
    .Q(\decoded_imm[1] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 _42242_ (.D(_02739_),
    .Q(\irq_pending[31] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _42243_ (.D(_02740_),
    .Q(\irq_pending[30] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 _42244_ (.D(_02741_),
    .Q(\irq_pending[29] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _42245_ (.D(_02742_),
    .Q(\irq_pending[28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_2 _42246_ (.D(_02743_),
    .Q(\irq_pending[27] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_2 _42247_ (.D(_02744_),
    .Q(\irq_pending[26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_2 _42248_ (.D(_02745_),
    .Q(\irq_pending[25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _42249_ (.D(_02746_),
    .Q(\irq_pending[24] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _42250_ (.D(_02747_),
    .Q(\irq_pending[23] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_1 _42251_ (.D(_02748_),
    .Q(\irq_pending[22] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_2 _42252_ (.D(_02749_),
    .Q(\irq_pending[21] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _42253_ (.D(_02750_),
    .Q(\irq_pending[20] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _42254_ (.D(_02751_),
    .Q(\irq_pending[19] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42255_ (.D(_02752_),
    .Q(\irq_pending[18] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _42256_ (.D(_02753_),
    .Q(\irq_pending[17] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_2 _42257_ (.D(_02754_),
    .Q(\irq_pending[16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_2 _42258_ (.D(_02755_),
    .Q(\irq_pending[15] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _42259_ (.D(_02756_),
    .Q(\irq_pending[14] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _42260_ (.D(_02757_),
    .Q(\irq_pending[13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _42261_ (.D(_02758_),
    .Q(\irq_pending[12] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _42262_ (.D(_02759_),
    .Q(\irq_pending[11] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_2 _42263_ (.D(_02760_),
    .Q(\irq_pending[10] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _42264_ (.D(_02761_),
    .Q(\irq_pending[9] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_2 _42265_ (.D(_02762_),
    .Q(\irq_pending[8] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _42266_ (.D(_02763_),
    .Q(\irq_pending[7] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _42267_ (.D(_02764_),
    .Q(\irq_pending[6] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _42268_ (.D(_02765_),
    .Q(\irq_pending[5] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _42269_ (.D(_02766_),
    .Q(\irq_pending[4] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_2 _42270_ (.D(_02767_),
    .Q(\irq_pending[3] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _42271_ (.D(_02768_),
    .Q(\irq_pending[1] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_2 _42272_ (.D(_02769_),
    .Q(\irq_pending[0] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_2 _42273_ (.D(_02770_),
    .Q(\reg_next_pc[0] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 _42274_ (.D(_00045_),
    .Q(\mem_wordsize[0] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_4 _42275_ (.D(_00046_),
    .Q(\mem_wordsize[1] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _42276_ (.D(_00047_),
    .Q(\mem_wordsize[2] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _42277_ (.D(_20896_),
    .Q(\reg_out[0] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _42278_ (.D(_20907_),
    .Q(\reg_out[1] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _42279_ (.D(_20918_),
    .Q(\reg_out[2] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 _42280_ (.D(_20921_),
    .Q(\reg_out[3] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 _42281_ (.D(_20922_),
    .Q(\reg_out[4] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 _42282_ (.D(_20923_),
    .Q(\reg_out[5] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 _42283_ (.D(_20924_),
    .Q(\reg_out[6] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 _42284_ (.D(_20925_),
    .Q(\reg_out[7] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__dfxtp_1 _42285_ (.D(_20926_),
    .Q(\reg_out[8] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 _42286_ (.D(_20927_),
    .Q(\reg_out[9] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _42287_ (.D(_20897_),
    .Q(\reg_out[10] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 _42288_ (.D(_20898_),
    .Q(\reg_out[11] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_1 _42289_ (.D(_20899_),
    .Q(\reg_out[12] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_1 _42290_ (.D(_20900_),
    .Q(\reg_out[13] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_1 _42291_ (.D(_20901_),
    .Q(\reg_out[14] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _42292_ (.D(_20902_),
    .Q(\reg_out[15] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _42293_ (.D(_20903_),
    .Q(\reg_out[16] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _42294_ (.D(_20904_),
    .Q(\reg_out[17] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _42295_ (.D(_20905_),
    .Q(\reg_out[18] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _42296_ (.D(_20906_),
    .Q(\reg_out[19] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _42297_ (.D(_20908_),
    .Q(\reg_out[20] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _42298_ (.D(_20909_),
    .Q(\reg_out[21] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _42299_ (.D(_20910_),
    .Q(\reg_out[22] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _42300_ (.D(_20911_),
    .Q(\reg_out[23] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_1 _42301_ (.D(_20912_),
    .Q(\reg_out[24] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _42302_ (.D(_20913_),
    .Q(\reg_out[25] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _42303_ (.D(_20914_),
    .Q(\reg_out[26] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__dfxtp_1 _42304_ (.D(_20915_),
    .Q(\reg_out[27] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 _42305_ (.D(_20916_),
    .Q(\reg_out[28] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 _42306_ (.D(_20917_),
    .Q(\reg_out[29] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _42307_ (.D(_20919_),
    .Q(\reg_out[30] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 _42308_ (.D(_20920_),
    .Q(\reg_out[31] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_2 _42309_ (.D(_00004_),
    .Q(\irq_pending[2] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_4 _42310_ (.D(_00003_),
    .Q(decoder_trigger),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_2 _42311_ (.D(\alu_out[0] ),
    .Q(\alu_out_q[0] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _42312_ (.D(\alu_out[1] ),
    .Q(\alu_out_q[1] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_2 _42313_ (.D(\alu_out[2] ),
    .Q(\alu_out_q[2] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_2 _42314_ (.D(\alu_out[3] ),
    .Q(\alu_out_q[3] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_2 _42315_ (.D(\alu_out[4] ),
    .Q(\alu_out_q[4] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 _42316_ (.D(\alu_out[5] ),
    .Q(\alu_out_q[5] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _42317_ (.D(\alu_out[6] ),
    .Q(\alu_out_q[6] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _42318_ (.D(\alu_out[7] ),
    .Q(\alu_out_q[7] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _42319_ (.D(\alu_out[8] ),
    .Q(\alu_out_q[8] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _42320_ (.D(\alu_out[9] ),
    .Q(\alu_out_q[9] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42321_ (.D(\alu_out[10] ),
    .Q(\alu_out_q[10] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _42322_ (.D(\alu_out[11] ),
    .Q(\alu_out_q[11] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42323_ (.D(\alu_out[12] ),
    .Q(\alu_out_q[12] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _42324_ (.D(\alu_out[13] ),
    .Q(\alu_out_q[13] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _42325_ (.D(\alu_out[14] ),
    .Q(\alu_out_q[14] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42326_ (.D(\alu_out[15] ),
    .Q(\alu_out_q[15] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42327_ (.D(\alu_out[16] ),
    .Q(\alu_out_q[16] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_1 _42328_ (.D(\alu_out[17] ),
    .Q(\alu_out_q[17] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42329_ (.D(\alu_out[18] ),
    .Q(\alu_out_q[18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_1 _42330_ (.D(\alu_out[19] ),
    .Q(\alu_out_q[19] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42331_ (.D(\alu_out[20] ),
    .Q(\alu_out_q[20] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _42332_ (.D(\alu_out[21] ),
    .Q(\alu_out_q[21] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_1 _42333_ (.D(\alu_out[22] ),
    .Q(\alu_out_q[22] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_1 _42334_ (.D(\alu_out[23] ),
    .Q(\alu_out_q[23] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_1 _42335_ (.D(\alu_out[24] ),
    .Q(\alu_out_q[24] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _42336_ (.D(\alu_out[25] ),
    .Q(\alu_out_q[25] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_2 _42337_ (.D(\alu_out[26] ),
    .Q(\alu_out_q[26] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 _42338_ (.D(\alu_out[27] ),
    .Q(\alu_out_q[27] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_2 _42339_ (.D(\alu_out[28] ),
    .Q(\alu_out_q[28] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_2 _42340_ (.D(\alu_out[29] ),
    .Q(\alu_out_q[29] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _42341_ (.D(\alu_out[30] ),
    .Q(\alu_out_q[30] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_2 _42342_ (.D(\alu_out[31] ),
    .Q(\alu_out_q[31] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_4 _42343_ (.D(_00005_),
    .Q(is_lui_auipc_jal),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 _42344_ (.D(_00006_),
    .Q(is_slti_blt_slt),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _42345_ (.D(_00007_),
    .Q(is_sltiu_bltu_sltu),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _42346_ (.D(_02591_),
    .Q(\alu_add_sub[0] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 _42347_ (.D(_02602_),
    .Q(\alu_add_sub[1] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 _42348_ (.D(_02613_),
    .Q(\alu_add_sub[2] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 _42349_ (.D(_02616_),
    .Q(\alu_add_sub[3] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 _42350_ (.D(_02617_),
    .Q(\alu_add_sub[4] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 _42351_ (.D(_02618_),
    .Q(\alu_add_sub[5] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 _42352_ (.D(_02619_),
    .Q(\alu_add_sub[6] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _42353_ (.D(_02620_),
    .Q(\alu_add_sub[7] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _42354_ (.D(_02621_),
    .Q(\alu_add_sub[8] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _42355_ (.D(_02622_),
    .Q(\alu_add_sub[9] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 _42356_ (.D(_02592_),
    .Q(\alu_add_sub[10] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _42357_ (.D(_02593_),
    .Q(\alu_add_sub[11] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42358_ (.D(_02594_),
    .Q(\alu_add_sub[12] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _42359_ (.D(_02595_),
    .Q(\alu_add_sub[13] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _42360_ (.D(_02596_),
    .Q(\alu_add_sub[14] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _42361_ (.D(_02597_),
    .Q(\alu_add_sub[15] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 _42362_ (.D(_02598_),
    .Q(\alu_add_sub[16] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _42363_ (.D(_02599_),
    .Q(\alu_add_sub[17] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _42364_ (.D(_02600_),
    .Q(\alu_add_sub[18] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _42365_ (.D(_02601_),
    .Q(\alu_add_sub[19] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _42366_ (.D(_02603_),
    .Q(\alu_add_sub[20] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42367_ (.D(_02604_),
    .Q(\alu_add_sub[21] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_1 _42368_ (.D(_02605_),
    .Q(\alu_add_sub[22] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_1 _42369_ (.D(_02606_),
    .Q(\alu_add_sub[23] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 _42370_ (.D(_02607_),
    .Q(\alu_add_sub[24] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 _42371_ (.D(_02608_),
    .Q(\alu_add_sub[25] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_1 _42372_ (.D(_02609_),
    .Q(\alu_add_sub[26] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 _42373_ (.D(_02610_),
    .Q(\alu_add_sub[27] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 _42374_ (.D(_02611_),
    .Q(\alu_add_sub[28] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 _42375_ (.D(_02612_),
    .Q(\alu_add_sub[29] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 _42376_ (.D(_02614_),
    .Q(\alu_add_sub[30] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 _42377_ (.D(_02615_),
    .Q(\alu_add_sub[31] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 _42378_ (.D(_20931_),
    .Q(\alu_shl[16] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42379_ (.D(_20932_),
    .Q(\alu_shl[17] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42380_ (.D(_20933_),
    .Q(\alu_shl[18] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42381_ (.D(_20934_),
    .Q(\alu_shl[19] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42382_ (.D(_20935_),
    .Q(\alu_shl[20] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42383_ (.D(_20936_),
    .Q(\alu_shl[21] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42384_ (.D(_20937_),
    .Q(\alu_shl[22] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42385_ (.D(_20938_),
    .Q(\alu_shl[23] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__dfxtp_1 _42386_ (.D(_20939_),
    .Q(\alu_shl[24] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42387_ (.D(_20940_),
    .Q(\alu_shl[25] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42388_ (.D(_20941_),
    .Q(\alu_shl[26] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 _42389_ (.D(_20942_),
    .Q(\alu_shl[27] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 _42390_ (.D(_20943_),
    .Q(\alu_shl[28] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_1 _42391_ (.D(_20944_),
    .Q(\alu_shl[29] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42392_ (.D(_20945_),
    .Q(\alu_shl[30] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42393_ (.D(_20946_),
    .Q(\alu_shl[31] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 _42394_ (.D(_20947_),
    .Q(\alu_shr[0] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42395_ (.D(_20958_),
    .Q(\alu_shr[1] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _42396_ (.D(_20969_),
    .Q(\alu_shr[2] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42397_ (.D(_20972_),
    .Q(\alu_shr[3] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42398_ (.D(_20973_),
    .Q(\alu_shr[4] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42399_ (.D(_20974_),
    .Q(\alu_shr[5] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42400_ (.D(_20975_),
    .Q(\alu_shr[6] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _42401_ (.D(_20976_),
    .Q(\alu_shr[7] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _42402_ (.D(_20977_),
    .Q(\alu_shr[8] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42403_ (.D(_20978_),
    .Q(\alu_shr[9] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _42404_ (.D(_20948_),
    .Q(\alu_shr[10] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42405_ (.D(_20949_),
    .Q(\alu_shr[11] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42406_ (.D(_20950_),
    .Q(\alu_shr[12] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42407_ (.D(_20951_),
    .Q(\alu_shr[13] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42408_ (.D(_20952_),
    .Q(\alu_shr[14] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _42409_ (.D(_20953_),
    .Q(\alu_shr[15] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _42410_ (.D(_20954_),
    .Q(\alu_shr[16] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42411_ (.D(_20955_),
    .Q(\alu_shr[17] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _42412_ (.D(_20956_),
    .Q(\alu_shr[18] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42413_ (.D(_20957_),
    .Q(\alu_shr[19] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42414_ (.D(_20959_),
    .Q(\alu_shr[20] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42415_ (.D(_20960_),
    .Q(\alu_shr[21] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42416_ (.D(_20961_),
    .Q(\alu_shr[22] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _42417_ (.D(_20962_),
    .Q(\alu_shr[23] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 _42418_ (.D(_20963_),
    .Q(\alu_shr[24] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42419_ (.D(_20964_),
    .Q(\alu_shr[25] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 _42420_ (.D(_20965_),
    .Q(\alu_shr[26] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 _42421_ (.D(_20966_),
    .Q(\alu_shr[27] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 _42422_ (.D(_20967_),
    .Q(\alu_shr[28] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 _42423_ (.D(_20968_),
    .Q(\alu_shr[29] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_2 _42424_ (.D(_20970_),
    .Q(\alu_shr[30] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _42425_ (.D(_20971_),
    .Q(\alu_shr[31] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _42426_ (.D(_00000_),
    .Q(alu_eq),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_2 _42427_ (.D(_00002_),
    .Q(alu_ltu),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_2 _42428_ (.D(_00001_),
    .Q(alu_lts),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42429_ (.D(_02623_),
    .Q(\pcpi_mul.rd[0] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 _42430_ (.D(_02624_),
    .Q(\pcpi_mul.rd[1] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 _42431_ (.D(_02625_),
    .Q(\pcpi_mul.rd[2] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_1 _42432_ (.D(_02626_),
    .Q(\pcpi_mul.rd[3] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_1 _42433_ (.D(_02627_),
    .Q(\pcpi_mul.rd[4] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__dfxtp_1 _42434_ (.D(_02628_),
    .Q(\pcpi_mul.rd[5] ),
    .CLK(clknet_5_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42435_ (.D(_02683_),
    .Q(\pcpi_mul.rd[6] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42436_ (.D(_02684_),
    .Q(\pcpi_mul.rd[7] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42437_ (.D(_02685_),
    .Q(\pcpi_mul.rd[8] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42438_ (.D(_02686_),
    .Q(\pcpi_mul.rd[9] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42439_ (.D(_02629_),
    .Q(\pcpi_mul.rd[10] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42440_ (.D(_02630_),
    .Q(\pcpi_mul.rd[11] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_4 _42441_ (.D(_02631_),
    .Q(\pcpi_mul.rd[12] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_4 _42442_ (.D(_02632_),
    .Q(\pcpi_mul.rd[13] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_4 _42443_ (.D(_02633_),
    .Q(\pcpi_mul.rd[14] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_4 _42444_ (.D(_02634_),
    .Q(\pcpi_mul.rd[15] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 _42445_ (.D(_02635_),
    .Q(\pcpi_mul.rd[16] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42446_ (.D(_02636_),
    .Q(\pcpi_mul.rd[17] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42447_ (.D(_02637_),
    .Q(\pcpi_mul.rd[18] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_2 _42448_ (.D(_02638_),
    .Q(\pcpi_mul.rd[19] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 _42449_ (.D(_02639_),
    .Q(\pcpi_mul.rd[20] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _42450_ (.D(_02640_),
    .Q(\pcpi_mul.rd[21] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42451_ (.D(_02641_),
    .Q(\pcpi_mul.rd[22] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__dfxtp_4 _42452_ (.D(_02642_),
    .Q(\pcpi_mul.rd[23] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _42453_ (.D(_02643_),
    .Q(\pcpi_mul.rd[24] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _42454_ (.D(_02644_),
    .Q(\pcpi_mul.rd[25] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 _42455_ (.D(_02645_),
    .Q(\pcpi_mul.rd[26] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 _42456_ (.D(_02646_),
    .Q(\pcpi_mul.rd[27] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _42457_ (.D(_02647_),
    .Q(\pcpi_mul.rd[28] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 _42458_ (.D(_02648_),
    .Q(\pcpi_mul.rd[29] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _42459_ (.D(_02649_),
    .Q(\pcpi_mul.rd[30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 _42460_ (.D(_02650_),
    .Q(\pcpi_mul.rd[31] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _42461_ (.D(_02651_),
    .Q(\pcpi_mul.rd[32] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 _42462_ (.D(_02652_),
    .Q(\pcpi_mul.rd[33] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 _42463_ (.D(_02653_),
    .Q(\pcpi_mul.rd[34] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__dfxtp_1 _42464_ (.D(_02654_),
    .Q(\pcpi_mul.rd[35] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 _42465_ (.D(_02655_),
    .Q(\pcpi_mul.rd[36] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 _42466_ (.D(_02656_),
    .Q(\pcpi_mul.rd[37] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 _42467_ (.D(_02657_),
    .Q(\pcpi_mul.rd[38] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 _42468_ (.D(_02658_),
    .Q(\pcpi_mul.rd[39] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 _42469_ (.D(_02659_),
    .Q(\pcpi_mul.rd[40] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 _42470_ (.D(_02660_),
    .Q(\pcpi_mul.rd[41] ),
    .CLK(clknet_5_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42471_ (.D(_02661_),
    .Q(\pcpi_mul.rd[42] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 _42472_ (.D(_02662_),
    .Q(\pcpi_mul.rd[43] ),
    .CLK(clknet_5_12_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42473_ (.D(_02663_),
    .Q(\pcpi_mul.rd[44] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 _42474_ (.D(_02664_),
    .Q(\pcpi_mul.rd[45] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 _42475_ (.D(_02665_),
    .Q(\pcpi_mul.rd[46] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_2 _42476_ (.D(_02666_),
    .Q(\pcpi_mul.rd[47] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _42477_ (.D(_02667_),
    .Q(\pcpi_mul.rd[48] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _42478_ (.D(_02668_),
    .Q(\pcpi_mul.rd[49] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _42479_ (.D(_02669_),
    .Q(\pcpi_mul.rd[50] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _42480_ (.D(_02670_),
    .Q(\pcpi_mul.rd[51] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 _42481_ (.D(_02671_),
    .Q(\pcpi_mul.rd[52] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _42482_ (.D(_02672_),
    .Q(\pcpi_mul.rd[53] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_4 _42483_ (.D(_02673_),
    .Q(\pcpi_mul.rd[54] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_4 _42484_ (.D(_02674_),
    .Q(\pcpi_mul.rd[55] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__dfxtp_1 _42485_ (.D(_02675_),
    .Q(\pcpi_mul.rd[56] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 _42486_ (.D(_02676_),
    .Q(\pcpi_mul.rd[57] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _42487_ (.D(_02677_),
    .Q(\pcpi_mul.rd[58] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _42488_ (.D(_02678_),
    .Q(\pcpi_mul.rd[59] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 _42489_ (.D(_02679_),
    .Q(\pcpi_mul.rd[60] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 _42490_ (.D(_02680_),
    .Q(\pcpi_mul.rd[61] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 _42491_ (.D(_02681_),
    .Q(\pcpi_mul.rd[62] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _42492_ (.D(_02682_),
    .Q(\pcpi_mul.rd[63] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_2 _42493_ (.D(\pcpi_mul.instr_any_mulh ),
    .Q(\pcpi_mul.shift_out ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 _42494_ (.D(_00038_),
    .Q(\cpu_state[0] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_2 _42495_ (.D(_00039_),
    .Q(\cpu_state[1] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_4 _42496_ (.D(_00040_),
    .Q(\cpu_state[2] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_4 _42497_ (.D(_00041_),
    .Q(\cpu_state[3] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_4 _42498_ (.D(_00042_),
    .Q(\cpu_state[4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_2 _42499_ (.D(_00043_),
    .Q(\cpu_state[5] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _42500_ (.D(_00044_),
    .Q(\cpu_state[6] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _42501_ (.D(_02771_),
    .Q(\cpuregs[8][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _42502_ (.D(_02772_),
    .Q(\cpuregs[8][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42503_ (.D(_02773_),
    .Q(\cpuregs[8][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _42504_ (.D(_02774_),
    .Q(\cpuregs[8][3] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _42505_ (.D(_02775_),
    .Q(\cpuregs[8][4] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42506_ (.D(_02776_),
    .Q(\cpuregs[8][5] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _42507_ (.D(_02777_),
    .Q(\cpuregs[8][6] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _42508_ (.D(_02778_),
    .Q(\cpuregs[8][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _42509_ (.D(_02779_),
    .Q(\cpuregs[8][8] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _42510_ (.D(_02780_),
    .Q(\cpuregs[8][9] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _42511_ (.D(_02781_),
    .Q(\cpuregs[8][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _42512_ (.D(_02782_),
    .Q(\cpuregs[8][11] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 _42513_ (.D(_02783_),
    .Q(\cpuregs[8][12] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _42514_ (.D(_02784_),
    .Q(\cpuregs[8][13] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _42515_ (.D(_02785_),
    .Q(\cpuregs[8][14] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _42516_ (.D(_02786_),
    .Q(\cpuregs[8][15] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _42517_ (.D(_02787_),
    .Q(\cpuregs[8][16] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _42518_ (.D(_02788_),
    .Q(\cpuregs[8][17] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _42519_ (.D(_02789_),
    .Q(\cpuregs[8][18] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _42520_ (.D(_02790_),
    .Q(\cpuregs[8][19] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _42521_ (.D(_02791_),
    .Q(\cpuregs[8][20] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _42522_ (.D(_02792_),
    .Q(\cpuregs[8][21] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _42523_ (.D(_02793_),
    .Q(\cpuregs[8][22] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _42524_ (.D(_02794_),
    .Q(\cpuregs[8][23] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _42525_ (.D(_02795_),
    .Q(\cpuregs[8][24] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _42526_ (.D(_02796_),
    .Q(\cpuregs[8][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _42527_ (.D(_02797_),
    .Q(\cpuregs[8][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _42528_ (.D(_02798_),
    .Q(\cpuregs[8][27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _42529_ (.D(_02799_),
    .Q(\cpuregs[8][28] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _42530_ (.D(_02800_),
    .Q(\cpuregs[8][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _42531_ (.D(_02801_),
    .Q(\cpuregs[8][30] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _42532_ (.D(_02802_),
    .Q(\cpuregs[8][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _42533_ (.D(_02803_),
    .Q(\cpuregs[14][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _42534_ (.D(_02804_),
    .Q(\cpuregs[14][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42535_ (.D(_02805_),
    .Q(\cpuregs[14][2] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _42536_ (.D(_02806_),
    .Q(\cpuregs[14][3] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _42537_ (.D(_02807_),
    .Q(\cpuregs[14][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _42538_ (.D(_02808_),
    .Q(\cpuregs[14][5] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _42539_ (.D(_02809_),
    .Q(\cpuregs[14][6] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _42540_ (.D(_02810_),
    .Q(\cpuregs[14][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _42541_ (.D(_02811_),
    .Q(\cpuregs[14][8] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _42542_ (.D(_02812_),
    .Q(\cpuregs[14][9] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _42543_ (.D(_02813_),
    .Q(\cpuregs[14][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _42544_ (.D(_02814_),
    .Q(\cpuregs[14][11] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 _42545_ (.D(_02815_),
    .Q(\cpuregs[14][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _42546_ (.D(_02816_),
    .Q(\cpuregs[14][13] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _42547_ (.D(_02817_),
    .Q(\cpuregs[14][14] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _42548_ (.D(_02818_),
    .Q(\cpuregs[14][15] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _42549_ (.D(_02819_),
    .Q(\cpuregs[14][16] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _42550_ (.D(_02820_),
    .Q(\cpuregs[14][17] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _42551_ (.D(_02821_),
    .Q(\cpuregs[14][18] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _42552_ (.D(_02822_),
    .Q(\cpuregs[14][19] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _42553_ (.D(_02823_),
    .Q(\cpuregs[14][20] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _42554_ (.D(_02824_),
    .Q(\cpuregs[14][21] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _42555_ (.D(_02825_),
    .Q(\cpuregs[14][22] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _42556_ (.D(_02826_),
    .Q(\cpuregs[14][23] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _42557_ (.D(_02827_),
    .Q(\cpuregs[14][24] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _42558_ (.D(_02828_),
    .Q(\cpuregs[14][25] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _42559_ (.D(_02829_),
    .Q(\cpuregs[14][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _42560_ (.D(_02830_),
    .Q(\cpuregs[14][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _42561_ (.D(_02831_),
    .Q(\cpuregs[14][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _42562_ (.D(_02832_),
    .Q(\cpuregs[14][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _42563_ (.D(_02833_),
    .Q(\cpuregs[14][30] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _42564_ (.D(_02834_),
    .Q(\cpuregs[14][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _42565_ (.D(_02835_),
    .Q(\cpuregs[0][0] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _42566_ (.D(_02836_),
    .Q(\cpuregs[0][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42567_ (.D(_02837_),
    .Q(\cpuregs[0][2] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 _42568_ (.D(_02838_),
    .Q(\cpuregs[0][3] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42569_ (.D(_02839_),
    .Q(\cpuregs[0][4] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 _42570_ (.D(_02840_),
    .Q(\cpuregs[0][5] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 _42571_ (.D(_02841_),
    .Q(\cpuregs[0][6] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _42572_ (.D(_02842_),
    .Q(\cpuregs[0][7] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _42573_ (.D(_02843_),
    .Q(\cpuregs[0][8] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _42574_ (.D(_02844_),
    .Q(\cpuregs[0][9] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _42575_ (.D(_02845_),
    .Q(\cpuregs[0][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _42576_ (.D(_02846_),
    .Q(\cpuregs[0][11] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _42577_ (.D(_02847_),
    .Q(\cpuregs[0][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _42578_ (.D(_02848_),
    .Q(\cpuregs[0][13] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _42579_ (.D(_02849_),
    .Q(\cpuregs[0][14] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _42580_ (.D(_02850_),
    .Q(\cpuregs[0][15] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _42581_ (.D(_02851_),
    .Q(\cpuregs[0][16] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _42582_ (.D(_02852_),
    .Q(\cpuregs[0][17] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _42583_ (.D(_02853_),
    .Q(\cpuregs[0][18] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42584_ (.D(_02854_),
    .Q(\cpuregs[0][19] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 _42585_ (.D(_02855_),
    .Q(\cpuregs[0][20] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _42586_ (.D(_02856_),
    .Q(\cpuregs[0][21] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42587_ (.D(_02857_),
    .Q(\cpuregs[0][22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _42588_ (.D(_02858_),
    .Q(\cpuregs[0][23] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _42589_ (.D(_02859_),
    .Q(\cpuregs[0][24] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _42590_ (.D(_02860_),
    .Q(\cpuregs[0][25] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _42591_ (.D(_02861_),
    .Q(\cpuregs[0][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _42592_ (.D(_02862_),
    .Q(\cpuregs[0][27] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _42593_ (.D(_02863_),
    .Q(\cpuregs[0][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _42594_ (.D(_02864_),
    .Q(\cpuregs[0][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _42595_ (.D(_02865_),
    .Q(\cpuregs[0][30] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _42596_ (.D(_02866_),
    .Q(\cpuregs[0][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _42597_ (.D(_02867_),
    .Q(\cpuregs[10][0] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _42598_ (.D(_02868_),
    .Q(\cpuregs[10][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42599_ (.D(_02869_),
    .Q(\cpuregs[10][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _42600_ (.D(_02870_),
    .Q(\cpuregs[10][3] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 _42601_ (.D(_02871_),
    .Q(\cpuregs[10][4] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 _42602_ (.D(_02872_),
    .Q(\cpuregs[10][5] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _42603_ (.D(_02873_),
    .Q(\cpuregs[10][6] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _42604_ (.D(_02874_),
    .Q(\cpuregs[10][7] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _42605_ (.D(_02875_),
    .Q(\cpuregs[10][8] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _42606_ (.D(_02876_),
    .Q(\cpuregs[10][9] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _42607_ (.D(_02877_),
    .Q(\cpuregs[10][10] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 _42608_ (.D(_02878_),
    .Q(\cpuregs[10][11] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 _42609_ (.D(_02879_),
    .Q(\cpuregs[10][12] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _42610_ (.D(_02880_),
    .Q(\cpuregs[10][13] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _42611_ (.D(_02881_),
    .Q(\cpuregs[10][14] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _42612_ (.D(_02882_),
    .Q(\cpuregs[10][15] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _42613_ (.D(_02883_),
    .Q(\cpuregs[10][16] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _42614_ (.D(_02884_),
    .Q(\cpuregs[10][17] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _42615_ (.D(_02885_),
    .Q(\cpuregs[10][18] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _42616_ (.D(_02886_),
    .Q(\cpuregs[10][19] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _42617_ (.D(_02887_),
    .Q(\cpuregs[10][20] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _42618_ (.D(_02888_),
    .Q(\cpuregs[10][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _42619_ (.D(_02889_),
    .Q(\cpuregs[10][22] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _42620_ (.D(_02890_),
    .Q(\cpuregs[10][23] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _42621_ (.D(_02891_),
    .Q(\cpuregs[10][24] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _42622_ (.D(_02892_),
    .Q(\cpuregs[10][25] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _42623_ (.D(_02893_),
    .Q(\cpuregs[10][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _42624_ (.D(_02894_),
    .Q(\cpuregs[10][27] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _42625_ (.D(_02895_),
    .Q(\cpuregs[10][28] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _42626_ (.D(_02896_),
    .Q(\cpuregs[10][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _42627_ (.D(_02897_),
    .Q(\cpuregs[10][30] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _42628_ (.D(_02898_),
    .Q(\cpuregs[10][31] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _42629_ (.D(_02899_),
    .Q(\cpuregs[18][0] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_1 _42630_ (.D(_02900_),
    .Q(\cpuregs[18][1] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 _42631_ (.D(_02901_),
    .Q(\cpuregs[18][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42632_ (.D(_02902_),
    .Q(\cpuregs[18][3] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _42633_ (.D(_02903_),
    .Q(\cpuregs[18][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _42634_ (.D(_02904_),
    .Q(\cpuregs[18][5] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _42635_ (.D(_02905_),
    .Q(\cpuregs[18][6] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _42636_ (.D(_02906_),
    .Q(\cpuregs[18][7] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _42637_ (.D(_02907_),
    .Q(\cpuregs[18][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _42638_ (.D(_02908_),
    .Q(\cpuregs[18][9] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _42639_ (.D(_02909_),
    .Q(\cpuregs[18][10] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 _42640_ (.D(_02910_),
    .Q(\cpuregs[18][11] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 _42641_ (.D(_02911_),
    .Q(\cpuregs[18][12] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _42642_ (.D(_02912_),
    .Q(\cpuregs[18][13] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _42643_ (.D(_02913_),
    .Q(\cpuregs[18][14] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _42644_ (.D(_02914_),
    .Q(\cpuregs[18][15] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _42645_ (.D(_02915_),
    .Q(\cpuregs[18][16] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _42646_ (.D(_02916_),
    .Q(\cpuregs[18][17] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _42647_ (.D(_02917_),
    .Q(\cpuregs[18][18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42648_ (.D(_02918_),
    .Q(\cpuregs[18][19] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42649_ (.D(_02919_),
    .Q(\cpuregs[18][20] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _42650_ (.D(_02920_),
    .Q(\cpuregs[18][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _42651_ (.D(_02921_),
    .Q(\cpuregs[18][22] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_1 _42652_ (.D(_02922_),
    .Q(\cpuregs[18][23] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _42653_ (.D(_02923_),
    .Q(\cpuregs[18][24] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _42654_ (.D(_02924_),
    .Q(\cpuregs[18][25] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _42655_ (.D(_02925_),
    .Q(\cpuregs[18][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _42656_ (.D(_02926_),
    .Q(\cpuregs[18][27] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _42657_ (.D(_02927_),
    .Q(\cpuregs[18][28] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _42658_ (.D(_02928_),
    .Q(\cpuregs[18][29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _42659_ (.D(_02929_),
    .Q(\cpuregs[18][30] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _42660_ (.D(_02930_),
    .Q(\cpuregs[18][31] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _42661_ (.D(_02931_),
    .Q(\mem_rdata_q[0] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 _42662_ (.D(_02932_),
    .Q(\mem_rdata_q[1] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 _42663_ (.D(_02933_),
    .Q(\mem_rdata_q[2] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 _42664_ (.D(_02934_),
    .Q(\mem_rdata_q[3] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 _42665_ (.D(_02935_),
    .Q(\mem_rdata_q[4] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 _42666_ (.D(_02936_),
    .Q(\mem_rdata_q[5] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 _42667_ (.D(_02937_),
    .Q(\mem_rdata_q[6] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _42668_ (.D(_02938_),
    .Q(\mem_rdata_q[7] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_2 _42669_ (.D(_02939_),
    .Q(\mem_rdata_q[8] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _42670_ (.D(_02940_),
    .Q(\mem_rdata_q[9] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_2 _42671_ (.D(_02941_),
    .Q(\mem_rdata_q[10] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_2 _42672_ (.D(_02942_),
    .Q(\mem_rdata_q[11] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_2 _42673_ (.D(_02943_),
    .Q(\mem_rdata_q[12] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_4 _42674_ (.D(_02944_),
    .Q(\mem_rdata_q[13] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_2 _42675_ (.D(_02945_),
    .Q(\mem_rdata_q[14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_2 _42676_ (.D(_02946_),
    .Q(\mem_rdata_q[15] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _42677_ (.D(_02947_),
    .Q(\mem_rdata_q[16] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_2 _42678_ (.D(_02948_),
    .Q(\mem_rdata_q[17] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_2 _42679_ (.D(_02949_),
    .Q(\mem_rdata_q[18] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_2 _42680_ (.D(_02950_),
    .Q(\mem_rdata_q[19] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 _42681_ (.D(_02951_),
    .Q(\mem_rdata_q[20] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 _42682_ (.D(_02952_),
    .Q(\mem_rdata_q[21] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_4 _42683_ (.D(_02953_),
    .Q(\mem_rdata_q[22] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42684_ (.D(_02954_),
    .Q(\mem_rdata_q[23] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_4 _42685_ (.D(_02955_),
    .Q(\mem_rdata_q[24] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_4 _42686_ (.D(_02956_),
    .Q(\mem_rdata_q[25] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _42687_ (.D(_02957_),
    .Q(\mem_rdata_q[26] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _42688_ (.D(_02958_),
    .Q(\mem_rdata_q[27] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42689_ (.D(_02959_),
    .Q(\mem_rdata_q[28] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42690_ (.D(_02960_),
    .Q(\mem_rdata_q[29] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _42691_ (.D(_02961_),
    .Q(\mem_rdata_q[30] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _42692_ (.D(_02962_),
    .Q(\mem_rdata_q[31] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 _42693_ (.D(_02963_),
    .Q(\cpuregs[2][0] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _42694_ (.D(_02964_),
    .Q(\cpuregs[2][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42695_ (.D(_02965_),
    .Q(\cpuregs[2][2] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 _42696_ (.D(_02966_),
    .Q(\cpuregs[2][3] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _42697_ (.D(_02967_),
    .Q(\cpuregs[2][4] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42698_ (.D(_02968_),
    .Q(\cpuregs[2][5] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 _42699_ (.D(_02969_),
    .Q(\cpuregs[2][6] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _42700_ (.D(_02970_),
    .Q(\cpuregs[2][7] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 _42701_ (.D(_02971_),
    .Q(\cpuregs[2][8] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _42702_ (.D(_02972_),
    .Q(\cpuregs[2][9] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _42703_ (.D(_02973_),
    .Q(\cpuregs[2][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _42704_ (.D(_02974_),
    .Q(\cpuregs[2][11] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _42705_ (.D(_02975_),
    .Q(\cpuregs[2][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _42706_ (.D(_02976_),
    .Q(\cpuregs[2][13] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _42707_ (.D(_02977_),
    .Q(\cpuregs[2][14] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _42708_ (.D(_02978_),
    .Q(\cpuregs[2][15] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _42709_ (.D(_02979_),
    .Q(\cpuregs[2][16] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _42710_ (.D(_02980_),
    .Q(\cpuregs[2][17] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _42711_ (.D(_02981_),
    .Q(\cpuregs[2][18] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _42712_ (.D(_02982_),
    .Q(\cpuregs[2][19] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _42713_ (.D(_02983_),
    .Q(\cpuregs[2][20] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _42714_ (.D(_02984_),
    .Q(\cpuregs[2][21] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _42715_ (.D(_02985_),
    .Q(\cpuregs[2][22] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42716_ (.D(_02986_),
    .Q(\cpuregs[2][23] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _42717_ (.D(_02987_),
    .Q(\cpuregs[2][24] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _42718_ (.D(_02988_),
    .Q(\cpuregs[2][25] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _42719_ (.D(_02989_),
    .Q(\cpuregs[2][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _42720_ (.D(_02990_),
    .Q(\cpuregs[2][27] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _42721_ (.D(_02991_),
    .Q(\cpuregs[2][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _42722_ (.D(_02992_),
    .Q(\cpuregs[2][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _42723_ (.D(_02993_),
    .Q(\cpuregs[2][30] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _42724_ (.D(_02994_),
    .Q(\cpuregs[2][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _42725_ (.D(_02995_),
    .Q(\cpuregs[5][0] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_1 _42726_ (.D(_02996_),
    .Q(\cpuregs[5][1] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _42727_ (.D(_02997_),
    .Q(\cpuregs[5][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _42728_ (.D(_02998_),
    .Q(\cpuregs[5][3] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _42729_ (.D(_02999_),
    .Q(\cpuregs[5][4] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _42730_ (.D(_03000_),
    .Q(\cpuregs[5][5] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _42731_ (.D(_03001_),
    .Q(\cpuregs[5][6] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _42732_ (.D(_03002_),
    .Q(\cpuregs[5][7] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _42733_ (.D(_03003_),
    .Q(\cpuregs[5][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _42734_ (.D(_03004_),
    .Q(\cpuregs[5][9] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _42735_ (.D(_03005_),
    .Q(\cpuregs[5][10] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 _42736_ (.D(_03006_),
    .Q(\cpuregs[5][11] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 _42737_ (.D(_03007_),
    .Q(\cpuregs[5][12] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _42738_ (.D(_03008_),
    .Q(\cpuregs[5][13] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _42739_ (.D(_03009_),
    .Q(\cpuregs[5][14] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _42740_ (.D(_03010_),
    .Q(\cpuregs[5][15] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _42741_ (.D(_03011_),
    .Q(\cpuregs[5][16] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _42742_ (.D(_03012_),
    .Q(\cpuregs[5][17] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _42743_ (.D(_03013_),
    .Q(\cpuregs[5][18] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _42744_ (.D(_03014_),
    .Q(\cpuregs[5][19] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _42745_ (.D(_03015_),
    .Q(\cpuregs[5][20] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _42746_ (.D(_03016_),
    .Q(\cpuregs[5][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _42747_ (.D(_03017_),
    .Q(\cpuregs[5][22] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_1 _42748_ (.D(_03018_),
    .Q(\cpuregs[5][23] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _42749_ (.D(_03019_),
    .Q(\cpuregs[5][24] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _42750_ (.D(_03020_),
    .Q(\cpuregs[5][25] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _42751_ (.D(_03021_),
    .Q(\cpuregs[5][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _42752_ (.D(_03022_),
    .Q(\cpuregs[5][27] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _42753_ (.D(_03023_),
    .Q(\cpuregs[5][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _42754_ (.D(_03024_),
    .Q(\cpuregs[5][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _42755_ (.D(_03025_),
    .Q(\cpuregs[5][30] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _42756_ (.D(_03026_),
    .Q(\cpuregs[5][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_4 _42757_ (.D(_03027_),
    .Q(\pcpi_mul.rs1[0] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 _42758_ (.D(_03028_),
    .Q(\pcpi_mul.rs1[1] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 _42759_ (.D(_03029_),
    .Q(\pcpi_mul.rs1[2] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 _42760_ (.D(_03030_),
    .Q(\pcpi_mul.rs1[3] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 _42761_ (.D(_03031_),
    .Q(\pcpi_mul.rs1[4] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_4 _42762_ (.D(_03032_),
    .Q(\pcpi_mul.rs1[5] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 _42763_ (.D(_03033_),
    .Q(\pcpi_mul.rs1[6] ),
    .CLK(clknet_5_13_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42764_ (.D(_03034_),
    .Q(\pcpi_mul.rs1[7] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 _42765_ (.D(_03035_),
    .Q(\pcpi_mul.rs1[8] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 _42766_ (.D(_03036_),
    .Q(\pcpi_mul.rs1[9] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 _42767_ (.D(_03037_),
    .Q(\pcpi_mul.rs1[10] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 _42768_ (.D(_03038_),
    .Q(\pcpi_mul.rs1[11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 _42769_ (.D(_03039_),
    .Q(\pcpi_mul.rs1[12] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_1 _42770_ (.D(_03040_),
    .Q(\pcpi_mul.rs1[13] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 _42771_ (.D(_03041_),
    .Q(\pcpi_mul.rs1[14] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _42772_ (.D(_03042_),
    .Q(\pcpi_mul.rs1[15] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _42773_ (.D(_03043_),
    .Q(\pcpi_mul.rs1[16] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _42774_ (.D(_03044_),
    .Q(\pcpi_mul.rs1[17] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__dfxtp_2 _42775_ (.D(_03045_),
    .Q(\pcpi_mul.rs1[18] ),
    .CLK(clknet_5_7_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42776_ (.D(_03046_),
    .Q(\pcpi_mul.rs1[19] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42777_ (.D(_03047_),
    .Q(\pcpi_mul.rs1[20] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_1 _42778_ (.D(_03048_),
    .Q(\pcpi_mul.rs1[21] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 _42779_ (.D(_03049_),
    .Q(\pcpi_mul.rs1[22] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_2 _42780_ (.D(_03050_),
    .Q(\pcpi_mul.rs1[23] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 _42781_ (.D(_03051_),
    .Q(\pcpi_mul.rs1[24] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42782_ (.D(_03052_),
    .Q(\pcpi_mul.rs1[25] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_1 _42783_ (.D(_03053_),
    .Q(\pcpi_mul.rs1[26] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_2 _42784_ (.D(_03054_),
    .Q(\pcpi_mul.rs1[27] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 _42785_ (.D(_03055_),
    .Q(\pcpi_mul.rs1[28] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_2 _42786_ (.D(_03056_),
    .Q(\pcpi_mul.rs1[29] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_4 _42787_ (.D(_03057_),
    .Q(\pcpi_mul.rs1[30] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_4 _42788_ (.D(_03058_),
    .Q(\pcpi_mul.rs1[31] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 _42789_ (.D(_03059_),
    .Q(net156),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_4 _42790_ (.D(_03060_),
    .Q(net159),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 _42791_ (.D(_03061_),
    .Q(net160),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _42792_ (.D(_03062_),
    .Q(net161),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_4 _42793_ (.D(_03063_),
    .Q(net162),
    .CLK(clknet_5_11_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _42794_ (.D(_03064_),
    .Q(net163),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _42795_ (.D(_03065_),
    .Q(net164),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 _42796_ (.D(_03066_),
    .Q(net165),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 _42797_ (.D(_03067_),
    .Q(net135),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _42798_ (.D(_03068_),
    .Q(net136),
    .CLK(clknet_5_10_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _42799_ (.D(_03069_),
    .Q(net137),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 _42800_ (.D(_03070_),
    .Q(net138),
    .CLK(clknet_5_15_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _42801_ (.D(_03071_),
    .Q(net139),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _42802_ (.D(_03072_),
    .Q(net140),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_2 _42803_ (.D(_03073_),
    .Q(net141),
    .CLK(clknet_5_31_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42804_ (.D(_03074_),
    .Q(net142),
    .CLK(clknet_opt_11_clk));
 sky130_fd_sc_hd__dfxtp_4 _42805_ (.D(_03075_),
    .Q(net143),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _42806_ (.D(_03076_),
    .Q(net144),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_4 _42807_ (.D(_03077_),
    .Q(net146),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _42808_ (.D(_03078_),
    .Q(net147),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 _42809_ (.D(_03079_),
    .Q(net148),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_4 _42810_ (.D(_03080_),
    .Q(net149),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_4 _42811_ (.D(_03081_),
    .Q(net150),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__dfxtp_4 _42812_ (.D(_03082_),
    .Q(net151),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_4 _42813_ (.D(_03083_),
    .Q(net152),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_4 _42814_ (.D(_03084_),
    .Q(net153),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _42815_ (.D(_03085_),
    .Q(net154),
    .CLK(clknet_5_10_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42816_ (.D(_03086_),
    .Q(net155),
    .CLK(clknet_5_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _42817_ (.D(_03087_),
    .Q(net157),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _42818_ (.D(_03088_),
    .Q(net158),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_4 _42819_ (.D(_03089_),
    .Q(net306),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _42820_ (.D(_03090_),
    .Q(net317),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_4 _42821_ (.D(_03091_),
    .Q(net328),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_4 _42822_ (.D(_03092_),
    .Q(net331),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_4 _42823_ (.D(_03093_),
    .Q(net332),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_4 _42824_ (.D(_03094_),
    .Q(net333),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_4 _42825_ (.D(_03095_),
    .Q(net334),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_4 _42826_ (.D(_03096_),
    .Q(net335),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_4 _42827_ (.D(_03097_),
    .Q(net336),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_4 _42828_ (.D(_03098_),
    .Q(net337),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__dfxtp_4 _42829_ (.D(_03099_),
    .Q(net307),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_4 _42830_ (.D(_03100_),
    .Q(net308),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_4 _42831_ (.D(_03101_),
    .Q(net309),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 _42832_ (.D(_03102_),
    .Q(net310),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 _42833_ (.D(_03103_),
    .Q(net311),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_4 _42834_ (.D(_03104_),
    .Q(net312),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_4 _42835_ (.D(_03105_),
    .Q(net313),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__dfxtp_4 _42836_ (.D(_03106_),
    .Q(net314),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_4 _42837_ (.D(_03107_),
    .Q(net315),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_4 _42838_ (.D(_03108_),
    .Q(net316),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_4 _42839_ (.D(_03109_),
    .Q(net318),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_4 _42840_ (.D(_03110_),
    .Q(net319),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_4 _42841_ (.D(_03111_),
    .Q(net320),
    .CLK(clknet_5_5_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _42842_ (.D(_03112_),
    .Q(net321),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_4 _42843_ (.D(_03113_),
    .Q(net322),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_4 _42844_ (.D(_03114_),
    .Q(net323),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_4 _42845_ (.D(_03115_),
    .Q(net324),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_4 _42846_ (.D(_03116_),
    .Q(net325),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_4 _42847_ (.D(_03117_),
    .Q(net326),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_4 _42848_ (.D(_03118_),
    .Q(net327),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_4 _42849_ (.D(_03119_),
    .Q(net329),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_4 _42850_ (.D(_03120_),
    .Q(net330),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_4 _42851_ (.D(_03121_),
    .Q(net274),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _42852_ (.D(_03122_),
    .Q(net285),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_4 _42853_ (.D(_03123_),
    .Q(net296),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _42854_ (.D(_03124_),
    .Q(net299),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42855_ (.D(_03125_),
    .Q(net300),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_4 _42856_ (.D(_03126_),
    .Q(net301),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _42857_ (.D(_03127_),
    .Q(net302),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42858_ (.D(_03128_),
    .Q(net303),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_2 _42859_ (.D(_03129_),
    .Q(net304),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42860_ (.D(_03130_),
    .Q(net305),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _42861_ (.D(_03131_),
    .Q(net275),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_4 _42862_ (.D(_03132_),
    .Q(net276),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_4 _42863_ (.D(_03133_),
    .Q(net277),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_4 _42864_ (.D(_03134_),
    .Q(net278),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _42865_ (.D(_03135_),
    .Q(net279),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _42866_ (.D(_03136_),
    .Q(net280),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_2 _42867_ (.D(_03137_),
    .Q(net281),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_4 _42868_ (.D(_03138_),
    .Q(net282),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _42869_ (.D(_03139_),
    .Q(net283),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _42870_ (.D(_03140_),
    .Q(net284),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_4 _42871_ (.D(_03141_),
    .Q(net286),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_4 _42872_ (.D(_03142_),
    .Q(net287),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42873_ (.D(_03143_),
    .Q(net288),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_4 _42874_ (.D(_03144_),
    .Q(net289),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_2 _42875_ (.D(_03145_),
    .Q(net290),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_4 _42876_ (.D(_03146_),
    .Q(net291),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_2 _42877_ (.D(_03147_),
    .Q(net292),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_4 _42878_ (.D(_03148_),
    .Q(net293),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_4 _42879_ (.D(_03149_),
    .Q(net294),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_4 _42880_ (.D(_03150_),
    .Q(net295),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_2 _42881_ (.D(_03151_),
    .Q(net297),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_4 _42882_ (.D(_03152_),
    .Q(net298),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_4 _42883_ (.D(_03153_),
    .Q(instr_lui),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_2 _42884_ (.D(_03154_),
    .Q(instr_auipc),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_4 _42885_ (.D(_03155_),
    .Q(instr_jal),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 _42886_ (.D(_03156_),
    .Q(instr_jalr),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 _42887_ (.D(_03157_),
    .Q(instr_lb),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _42888_ (.D(_03158_),
    .Q(instr_lh),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _42889_ (.D(_03159_),
    .Q(instr_lw),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _42890_ (.D(_03160_),
    .Q(instr_lbu),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _42891_ (.D(_03161_),
    .Q(instr_lhu),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _42892_ (.D(_03162_),
    .Q(instr_sb),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 _42893_ (.D(_03163_),
    .Q(instr_sh),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _42894_ (.D(_03164_),
    .Q(instr_sw),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _42895_ (.D(_03165_),
    .Q(instr_slli),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _42896_ (.D(_03166_),
    .Q(instr_srli),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 _42897_ (.D(_03167_),
    .Q(instr_srai),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 _42898_ (.D(_03168_),
    .Q(instr_rdcycle),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_2 _42899_ (.D(_03169_),
    .Q(instr_rdcycleh),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 _42900_ (.D(_03170_),
    .Q(instr_rdinstr),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_2 _42901_ (.D(_03171_),
    .Q(instr_rdinstrh),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_2 _42902_ (.D(_03172_),
    .Q(instr_ecall_ebreak),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _42903_ (.D(_03173_),
    .Q(instr_getq),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_2 _42904_ (.D(_03174_),
    .Q(instr_setq),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _42905_ (.D(_03175_),
    .Q(instr_retirq),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _42906_ (.D(_03176_),
    .Q(instr_maskirq),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_2 _42907_ (.D(_03177_),
    .Q(instr_waitirq),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_4 _42908_ (.D(_03178_),
    .Q(instr_timer),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfxtp_1 _42909_ (.D(_03179_),
    .Q(\decoded_rd[0] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_4 _42910_ (.D(_03180_),
    .Q(\decoded_rd[1] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_4 _42911_ (.D(_03181_),
    .Q(\decoded_rd[2] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_4 _42912_ (.D(_03182_),
    .Q(\decoded_rd[3] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _42913_ (.D(_03183_),
    .Q(\decoded_rd[4] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_2 _42914_ (.D(_03184_),
    .Q(\decoded_imm[0] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_4 _42915_ (.D(_03185_),
    .Q(\decoded_imm_uj[1] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_2 _42916_ (.D(_03186_),
    .Q(\decoded_imm_uj[2] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_4 _42917_ (.D(_03187_),
    .Q(\decoded_imm_uj[3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_4 _42918_ (.D(_03188_),
    .Q(\decoded_imm_uj[4] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42919_ (.D(_03189_),
    .Q(\decoded_imm_uj[5] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_2 _42920_ (.D(_03190_),
    .Q(\decoded_imm_uj[6] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_4 _42921_ (.D(_03191_),
    .Q(\decoded_imm_uj[7] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 _42922_ (.D(_03192_),
    .Q(\decoded_imm_uj[8] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_2 _42923_ (.D(_03193_),
    .Q(\decoded_imm_uj[9] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _42924_ (.D(_03194_),
    .Q(\decoded_imm_uj[10] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _42925_ (.D(_03195_),
    .Q(\decoded_imm_uj[11] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_4 _42926_ (.D(_03196_),
    .Q(\decoded_imm_uj[12] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_4 _42927_ (.D(_03197_),
    .Q(\decoded_imm_uj[13] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_4 _42928_ (.D(_03198_),
    .Q(\decoded_imm_uj[14] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_2 _42929_ (.D(_03199_),
    .Q(\decoded_imm_uj[15] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_2 _42930_ (.D(_03200_),
    .Q(\decoded_imm_uj[16] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_2 _42931_ (.D(_03201_),
    .Q(\decoded_imm_uj[17] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_2 _42932_ (.D(_03202_),
    .Q(\decoded_imm_uj[18] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_4 _42933_ (.D(_03203_),
    .Q(\decoded_imm_uj[19] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 _42934_ (.D(_03204_),
    .Q(\decoded_imm_uj[20] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _42935_ (.D(_03205_),
    .Q(is_lb_lh_lw_lbu_lhu),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_4 _42936_ (.D(_03206_),
    .Q(is_slli_srli_srai),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_4 _42937_ (.D(_03207_),
    .Q(is_jalr_addi_slti_sltiu_xori_ori_andi),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_2 _42938_ (.D(_03208_),
    .Q(is_sb_sh_sw),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 _42939_ (.D(_03209_),
    .Q(\cpuregs[13][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _42940_ (.D(_03210_),
    .Q(\cpuregs[13][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _42941_ (.D(_03211_),
    .Q(\cpuregs[13][2] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _42942_ (.D(_03212_),
    .Q(\cpuregs[13][3] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _42943_ (.D(_03213_),
    .Q(\cpuregs[13][4] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _42944_ (.D(_03214_),
    .Q(\cpuregs[13][5] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _42945_ (.D(_03215_),
    .Q(\cpuregs[13][6] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _42946_ (.D(_03216_),
    .Q(\cpuregs[13][7] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _42947_ (.D(_03217_),
    .Q(\cpuregs[13][8] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _42948_ (.D(_03218_),
    .Q(\cpuregs[13][9] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _42949_ (.D(_03219_),
    .Q(\cpuregs[13][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _42950_ (.D(_03220_),
    .Q(\cpuregs[13][11] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _42951_ (.D(_03221_),
    .Q(\cpuregs[13][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _42952_ (.D(_03222_),
    .Q(\cpuregs[13][13] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _42953_ (.D(_03223_),
    .Q(\cpuregs[13][14] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _42954_ (.D(_03224_),
    .Q(\cpuregs[13][15] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _42955_ (.D(_03225_),
    .Q(\cpuregs[13][16] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _42956_ (.D(_03226_),
    .Q(\cpuregs[13][17] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _42957_ (.D(_03227_),
    .Q(\cpuregs[13][18] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _42958_ (.D(_03228_),
    .Q(\cpuregs[13][19] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 _42959_ (.D(_03229_),
    .Q(\cpuregs[13][20] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _42960_ (.D(_03230_),
    .Q(\cpuregs[13][21] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _42961_ (.D(_03231_),
    .Q(\cpuregs[13][22] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _42962_ (.D(_03232_),
    .Q(\cpuregs[13][23] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _42963_ (.D(_03233_),
    .Q(\cpuregs[13][24] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _42964_ (.D(_03234_),
    .Q(\cpuregs[13][25] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _42965_ (.D(_03235_),
    .Q(\cpuregs[13][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _42966_ (.D(_03236_),
    .Q(\cpuregs[13][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _42967_ (.D(_03237_),
    .Q(\cpuregs[13][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _42968_ (.D(_03238_),
    .Q(\cpuregs[13][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _42969_ (.D(_03239_),
    .Q(\cpuregs[13][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _42970_ (.D(_03240_),
    .Q(\cpuregs[13][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _42971_ (.D(_03241_),
    .Q(is_alu_reg_imm),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 _42972_ (.D(_03242_),
    .Q(is_alu_reg_reg),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_4 _42973_ (.D(_03243_),
    .Q(net270),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_4 _42974_ (.D(_03244_),
    .Q(net271),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_4 _42975_ (.D(_03245_),
    .Q(net272),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_4 _42976_ (.D(_03246_),
    .Q(net273),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_4 _42977_ (.D(_03247_),
    .Q(\pcpi_mul.rs2[0] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__dfxtp_1 _42978_ (.D(_03248_),
    .Q(\pcpi_mul.rs2[1] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_1 _42979_ (.D(_03249_),
    .Q(\pcpi_mul.rs2[2] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_1 _42980_ (.D(_03250_),
    .Q(\pcpi_mul.rs2[3] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_2 _42981_ (.D(_03251_),
    .Q(\pcpi_mul.rs2[4] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__dfxtp_1 _42982_ (.D(_03252_),
    .Q(\pcpi_mul.rs2[5] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_4 _42983_ (.D(_03253_),
    .Q(\pcpi_mul.rs2[6] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 _42984_ (.D(_03254_),
    .Q(\pcpi_mul.rs2[7] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 _42985_ (.D(_03255_),
    .Q(\pcpi_mul.rs2[8] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__dfxtp_1 _42986_ (.D(_03256_),
    .Q(\pcpi_mul.rs2[9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _42987_ (.D(_03257_),
    .Q(\pcpi_mul.rs2[10] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _42988_ (.D(_03258_),
    .Q(\pcpi_mul.rs2[11] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_4 _42989_ (.D(_03259_),
    .Q(\pcpi_mul.rs2[12] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__dfxtp_1 _42990_ (.D(_03260_),
    .Q(\pcpi_mul.rs2[13] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_1 _42991_ (.D(_03261_),
    .Q(\pcpi_mul.rs2[14] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__dfxtp_2 _42992_ (.D(_03262_),
    .Q(\pcpi_mul.rs2[15] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 _42993_ (.D(_03263_),
    .Q(\pcpi_mul.rs2[16] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__dfxtp_2 _42994_ (.D(_03264_),
    .Q(\pcpi_mul.rs2[17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_4 _42995_ (.D(_03265_),
    .Q(\pcpi_mul.rs2[18] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_1 _42996_ (.D(_03266_),
    .Q(\pcpi_mul.rs2[19] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_2 _42997_ (.D(_03267_),
    .Q(\pcpi_mul.rs2[20] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dfxtp_2 _42998_ (.D(_03268_),
    .Q(\pcpi_mul.rs2[21] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_2 _42999_ (.D(_03269_),
    .Q(\pcpi_mul.rs2[22] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_2 _43000_ (.D(_03270_),
    .Q(\pcpi_mul.rs2[23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_4 _43001_ (.D(_03271_),
    .Q(\pcpi_mul.rs2[24] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_2 _43002_ (.D(_03272_),
    .Q(\pcpi_mul.rs2[25] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__dfxtp_4 _43003_ (.D(_03273_),
    .Q(\pcpi_mul.rs2[26] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__dfxtp_4 _43004_ (.D(_03274_),
    .Q(\pcpi_mul.rs2[27] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_4 _43005_ (.D(_03275_),
    .Q(\pcpi_mul.rs2[28] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__dfxtp_4 _43006_ (.D(_03276_),
    .Q(\pcpi_mul.rs2[29] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_4 _43007_ (.D(_03277_),
    .Q(\pcpi_mul.rs2[30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_4 _43008_ (.D(_03278_),
    .Q(\pcpi_mul.rs2[31] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _43009_ (.D(_03279_),
    .Q(\cpuregs[17][0] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _43010_ (.D(_03280_),
    .Q(\cpuregs[17][1] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_1 _43011_ (.D(_03281_),
    .Q(\cpuregs[17][2] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _43012_ (.D(_03282_),
    .Q(\cpuregs[17][3] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43013_ (.D(_03283_),
    .Q(\cpuregs[17][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43014_ (.D(_03284_),
    .Q(\cpuregs[17][5] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43015_ (.D(_03285_),
    .Q(\cpuregs[17][6] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43016_ (.D(_03286_),
    .Q(\cpuregs[17][7] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43017_ (.D(_03287_),
    .Q(\cpuregs[17][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _43018_ (.D(_03288_),
    .Q(\cpuregs[17][9] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43019_ (.D(_03289_),
    .Q(\cpuregs[17][10] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _43020_ (.D(_03290_),
    .Q(\cpuregs[17][11] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 _43021_ (.D(_03291_),
    .Q(\cpuregs[17][12] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43022_ (.D(_03292_),
    .Q(\cpuregs[17][13] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43023_ (.D(_03293_),
    .Q(\cpuregs[17][14] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43024_ (.D(_03294_),
    .Q(\cpuregs[17][15] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43025_ (.D(_03295_),
    .Q(\cpuregs[17][16] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _43026_ (.D(_03296_),
    .Q(\cpuregs[17][17] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43027_ (.D(_03297_),
    .Q(\cpuregs[17][18] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _43028_ (.D(_03298_),
    .Q(\cpuregs[17][19] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _43029_ (.D(_03299_),
    .Q(\cpuregs[17][20] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _43030_ (.D(_03300_),
    .Q(\cpuregs[17][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43031_ (.D(_03301_),
    .Q(\cpuregs[17][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _43032_ (.D(_03302_),
    .Q(\cpuregs[17][23] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _43033_ (.D(_03303_),
    .Q(\cpuregs[17][24] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43034_ (.D(_03304_),
    .Q(\cpuregs[17][25] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _43035_ (.D(_03305_),
    .Q(\cpuregs[17][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43036_ (.D(_03306_),
    .Q(\cpuregs[17][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43037_ (.D(_03307_),
    .Q(\cpuregs[17][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43038_ (.D(_03308_),
    .Q(\cpuregs[17][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _43039_ (.D(_03309_),
    .Q(\cpuregs[17][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43040_ (.D(_03310_),
    .Q(\cpuregs[17][31] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43041_ (.D(_03311_),
    .Q(\cpuregs[16][0] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _43042_ (.D(_03312_),
    .Q(\cpuregs[16][1] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_1 _43043_ (.D(_03313_),
    .Q(\cpuregs[16][2] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _43044_ (.D(_03314_),
    .Q(\cpuregs[16][3] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43045_ (.D(_03315_),
    .Q(\cpuregs[16][4] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 _43046_ (.D(_03316_),
    .Q(\cpuregs[16][5] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43047_ (.D(_03317_),
    .Q(\cpuregs[16][6] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43048_ (.D(_03318_),
    .Q(\cpuregs[16][7] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43049_ (.D(_03319_),
    .Q(\cpuregs[16][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _43050_ (.D(_03320_),
    .Q(\cpuregs[16][9] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43051_ (.D(_03321_),
    .Q(\cpuregs[16][10] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _43052_ (.D(_03322_),
    .Q(\cpuregs[16][11] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _43053_ (.D(_03323_),
    .Q(\cpuregs[16][12] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43054_ (.D(_03324_),
    .Q(\cpuregs[16][13] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43055_ (.D(_03325_),
    .Q(\cpuregs[16][14] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43056_ (.D(_03326_),
    .Q(\cpuregs[16][15] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43057_ (.D(_03327_),
    .Q(\cpuregs[16][16] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43058_ (.D(_03328_),
    .Q(\cpuregs[16][17] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43059_ (.D(_03329_),
    .Q(\cpuregs[16][18] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 _43060_ (.D(_03330_),
    .Q(\cpuregs[16][19] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 _43061_ (.D(_03331_),
    .Q(\cpuregs[16][20] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43062_ (.D(_03332_),
    .Q(\cpuregs[16][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43063_ (.D(_03333_),
    .Q(\cpuregs[16][22] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43064_ (.D(_03334_),
    .Q(\cpuregs[16][23] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _43065_ (.D(_03335_),
    .Q(\cpuregs[16][24] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43066_ (.D(_03336_),
    .Q(\cpuregs[16][25] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _43067_ (.D(_03337_),
    .Q(\cpuregs[16][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43068_ (.D(_03338_),
    .Q(\cpuregs[16][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43069_ (.D(_03339_),
    .Q(\cpuregs[16][28] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _43070_ (.D(_03340_),
    .Q(\cpuregs[16][29] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43071_ (.D(_03341_),
    .Q(\cpuregs[16][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43072_ (.D(_03342_),
    .Q(\cpuregs[16][31] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43073_ (.D(_03343_),
    .Q(\cpuregs[12][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _43074_ (.D(_03344_),
    .Q(\cpuregs[12][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _43075_ (.D(_03345_),
    .Q(\cpuregs[12][2] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _43076_ (.D(_03346_),
    .Q(\cpuregs[12][3] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43077_ (.D(_03347_),
    .Q(\cpuregs[12][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43078_ (.D(_03348_),
    .Q(\cpuregs[12][5] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _43079_ (.D(_03349_),
    .Q(\cpuregs[12][6] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 _43080_ (.D(_03350_),
    .Q(\cpuregs[12][7] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _43081_ (.D(_03351_),
    .Q(\cpuregs[12][8] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _43082_ (.D(_03352_),
    .Q(\cpuregs[12][9] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43083_ (.D(_03353_),
    .Q(\cpuregs[12][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43084_ (.D(_03354_),
    .Q(\cpuregs[12][11] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _43085_ (.D(_03355_),
    .Q(\cpuregs[12][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43086_ (.D(_03356_),
    .Q(\cpuregs[12][13] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43087_ (.D(_03357_),
    .Q(\cpuregs[12][14] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43088_ (.D(_03358_),
    .Q(\cpuregs[12][15] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43089_ (.D(_03359_),
    .Q(\cpuregs[12][16] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43090_ (.D(_03360_),
    .Q(\cpuregs[12][17] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43091_ (.D(_03361_),
    .Q(\cpuregs[12][18] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _43092_ (.D(_03362_),
    .Q(\cpuregs[12][19] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 _43093_ (.D(_03363_),
    .Q(\cpuregs[12][20] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43094_ (.D(_03364_),
    .Q(\cpuregs[12][21] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43095_ (.D(_03365_),
    .Q(\cpuregs[12][22] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43096_ (.D(_03366_),
    .Q(\cpuregs[12][23] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__dfxtp_1 _43097_ (.D(_03367_),
    .Q(\cpuregs[12][24] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43098_ (.D(_03368_),
    .Q(\cpuregs[12][25] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43099_ (.D(_03369_),
    .Q(\cpuregs[12][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _43100_ (.D(_03370_),
    .Q(\cpuregs[12][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43101_ (.D(_03371_),
    .Q(\cpuregs[12][28] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _43102_ (.D(_03372_),
    .Q(\cpuregs[12][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _43103_ (.D(_03373_),
    .Q(\cpuregs[12][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43104_ (.D(_03374_),
    .Q(\cpuregs[12][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43105_ (.D(_03375_),
    .Q(\cpuregs[1][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _43106_ (.D(_03376_),
    .Q(\cpuregs[1][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _43107_ (.D(_03377_),
    .Q(\cpuregs[1][2] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _43108_ (.D(_03378_),
    .Q(\cpuregs[1][3] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _43109_ (.D(_03379_),
    .Q(\cpuregs[1][4] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 _43110_ (.D(_03380_),
    .Q(\cpuregs[1][5] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _43111_ (.D(_03381_),
    .Q(\cpuregs[1][6] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _43112_ (.D(_03382_),
    .Q(\cpuregs[1][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _43113_ (.D(_03383_),
    .Q(\cpuregs[1][8] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _43114_ (.D(_03384_),
    .Q(\cpuregs[1][9] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _43115_ (.D(_03385_),
    .Q(\cpuregs[1][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _43116_ (.D(_03386_),
    .Q(\cpuregs[1][11] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _43117_ (.D(_03387_),
    .Q(\cpuregs[1][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _43118_ (.D(_03388_),
    .Q(\cpuregs[1][13] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43119_ (.D(_03389_),
    .Q(\cpuregs[1][14] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43120_ (.D(_03390_),
    .Q(\cpuregs[1][15] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43121_ (.D(_03391_),
    .Q(\cpuregs[1][16] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43122_ (.D(_03392_),
    .Q(\cpuregs[1][17] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__dfxtp_1 _43123_ (.D(_03393_),
    .Q(\cpuregs[1][18] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _43124_ (.D(_03394_),
    .Q(\cpuregs[1][19] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 _43125_ (.D(_03395_),
    .Q(\cpuregs[1][20] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _43126_ (.D(_03396_),
    .Q(\cpuregs[1][21] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43127_ (.D(_03397_),
    .Q(\cpuregs[1][22] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43128_ (.D(_03398_),
    .Q(\cpuregs[1][23] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _43129_ (.D(_03399_),
    .Q(\cpuregs[1][24] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43130_ (.D(_03400_),
    .Q(\cpuregs[1][25] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43131_ (.D(_03401_),
    .Q(\cpuregs[1][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43132_ (.D(_03402_),
    .Q(\cpuregs[1][27] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _43133_ (.D(_03403_),
    .Q(\cpuregs[1][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43134_ (.D(_03404_),
    .Q(\cpuregs[1][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _43135_ (.D(_03405_),
    .Q(\cpuregs[1][30] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _43136_ (.D(_03406_),
    .Q(\cpuregs[1][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43137_ (.D(_03407_),
    .Q(\cpuregs[3][0] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _43138_ (.D(_03408_),
    .Q(\cpuregs[3][1] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _43139_ (.D(_03409_),
    .Q(\cpuregs[3][2] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__dfxtp_1 _43140_ (.D(_03410_),
    .Q(\cpuregs[3][3] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _43141_ (.D(_03411_),
    .Q(\cpuregs[3][4] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 _43142_ (.D(_03412_),
    .Q(\cpuregs[3][5] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__dfxtp_1 _43143_ (.D(_03413_),
    .Q(\cpuregs[3][6] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _43144_ (.D(_03414_),
    .Q(\cpuregs[3][7] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _43145_ (.D(_03415_),
    .Q(\cpuregs[3][8] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _43146_ (.D(_03416_),
    .Q(\cpuregs[3][9] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 _43147_ (.D(_03417_),
    .Q(\cpuregs[3][10] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _43148_ (.D(_03418_),
    .Q(\cpuregs[3][11] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 _43149_ (.D(_03419_),
    .Q(\cpuregs[3][12] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 _43150_ (.D(_03420_),
    .Q(\cpuregs[3][13] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43151_ (.D(_03421_),
    .Q(\cpuregs[3][14] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 _43152_ (.D(_03422_),
    .Q(\cpuregs[3][15] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43153_ (.D(_03423_),
    .Q(\cpuregs[3][16] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_1 _43154_ (.D(_03424_),
    .Q(\cpuregs[3][17] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43155_ (.D(_03425_),
    .Q(\cpuregs[3][18] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _43156_ (.D(_03426_),
    .Q(\cpuregs[3][19] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _43157_ (.D(_03427_),
    .Q(\cpuregs[3][20] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43158_ (.D(_03428_),
    .Q(\cpuregs[3][21] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43159_ (.D(_03429_),
    .Q(\cpuregs[3][22] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43160_ (.D(_03430_),
    .Q(\cpuregs[3][23] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__dfxtp_1 _43161_ (.D(_03431_),
    .Q(\cpuregs[3][24] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43162_ (.D(_03432_),
    .Q(\cpuregs[3][25] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__dfxtp_1 _43163_ (.D(_03433_),
    .Q(\cpuregs[3][26] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 _43164_ (.D(_03434_),
    .Q(\cpuregs[3][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _43165_ (.D(_03435_),
    .Q(\cpuregs[3][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43166_ (.D(_03436_),
    .Q(\cpuregs[3][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _43167_ (.D(_03437_),
    .Q(\cpuregs[3][30] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _43168_ (.D(_03438_),
    .Q(\cpuregs[3][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 _43169_ (.D(_03439_),
    .Q(\cpuregs[11][0] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__dfxtp_1 _43170_ (.D(_03440_),
    .Q(\cpuregs[11][1] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _43171_ (.D(_03441_),
    .Q(\cpuregs[11][2] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _43172_ (.D(_03442_),
    .Q(\cpuregs[11][3] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _43173_ (.D(_03443_),
    .Q(\cpuregs[11][4] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _43174_ (.D(_03444_),
    .Q(\cpuregs[11][5] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 _43175_ (.D(_03445_),
    .Q(\cpuregs[11][6] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43176_ (.D(_03446_),
    .Q(\cpuregs[11][7] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _43177_ (.D(_03447_),
    .Q(\cpuregs[11][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _43178_ (.D(_03448_),
    .Q(\cpuregs[11][9] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _43179_ (.D(_03449_),
    .Q(\cpuregs[11][10] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 _43180_ (.D(_03450_),
    .Q(\cpuregs[11][11] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43181_ (.D(_03451_),
    .Q(\cpuregs[11][12] ),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfxtp_1 _43182_ (.D(_03452_),
    .Q(\cpuregs[11][13] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 _43183_ (.D(_03453_),
    .Q(\cpuregs[11][14] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43184_ (.D(_03454_),
    .Q(\cpuregs[11][15] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__dfxtp_1 _43185_ (.D(_03455_),
    .Q(\cpuregs[11][16] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _43186_ (.D(_03456_),
    .Q(\cpuregs[11][17] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 _43187_ (.D(_03457_),
    .Q(\cpuregs[11][18] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 _43188_ (.D(_03458_),
    .Q(\cpuregs[11][19] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _43189_ (.D(_03459_),
    .Q(\cpuregs[11][20] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43190_ (.D(_03460_),
    .Q(\cpuregs[11][21] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43191_ (.D(_03461_),
    .Q(\cpuregs[11][22] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43192_ (.D(_03462_),
    .Q(\cpuregs[11][23] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__dfxtp_1 _43193_ (.D(_03463_),
    .Q(\cpuregs[11][24] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43194_ (.D(_03464_),
    .Q(\cpuregs[11][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43195_ (.D(_03465_),
    .Q(\cpuregs[11][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43196_ (.D(_03466_),
    .Q(\cpuregs[11][27] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43197_ (.D(_03467_),
    .Q(\cpuregs[11][28] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 _43198_ (.D(_03468_),
    .Q(\cpuregs[11][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _43199_ (.D(_03469_),
    .Q(\cpuregs[11][30] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _43200_ (.D(_03470_),
    .Q(\cpuregs[11][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43201_ (.D(_03471_),
    .Q(\cpuregs[15][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _43202_ (.D(_03472_),
    .Q(\cpuregs[15][1] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 _43203_ (.D(_03473_),
    .Q(\cpuregs[15][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _43204_ (.D(_03474_),
    .Q(\cpuregs[15][3] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _43205_ (.D(_03475_),
    .Q(\cpuregs[15][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43206_ (.D(_03476_),
    .Q(\cpuregs[15][5] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__dfxtp_1 _43207_ (.D(_03477_),
    .Q(\cpuregs[15][6] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 _43208_ (.D(_03478_),
    .Q(\cpuregs[15][7] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _43209_ (.D(_03479_),
    .Q(\cpuregs[15][8] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 _43210_ (.D(_03480_),
    .Q(\cpuregs[15][9] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43211_ (.D(_03481_),
    .Q(\cpuregs[15][10] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43212_ (.D(_03482_),
    .Q(\cpuregs[15][11] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 _43213_ (.D(_03483_),
    .Q(\cpuregs[15][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43214_ (.D(_03484_),
    .Q(\cpuregs[15][13] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43215_ (.D(_03485_),
    .Q(\cpuregs[15][14] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43216_ (.D(_03486_),
    .Q(\cpuregs[15][15] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43217_ (.D(_03487_),
    .Q(\cpuregs[15][16] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43218_ (.D(_03488_),
    .Q(\cpuregs[15][17] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43219_ (.D(_03489_),
    .Q(\cpuregs[15][18] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _43220_ (.D(_03490_),
    .Q(\cpuregs[15][19] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _43221_ (.D(_03491_),
    .Q(\cpuregs[15][20] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43222_ (.D(_03492_),
    .Q(\cpuregs[15][21] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43223_ (.D(_03493_),
    .Q(\cpuregs[15][22] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43224_ (.D(_03494_),
    .Q(\cpuregs[15][23] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43225_ (.D(_03495_),
    .Q(\cpuregs[15][24] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43226_ (.D(_03496_),
    .Q(\cpuregs[15][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43227_ (.D(_03497_),
    .Q(\cpuregs[15][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _43228_ (.D(_03498_),
    .Q(\cpuregs[15][27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _43229_ (.D(_03499_),
    .Q(\cpuregs[15][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43230_ (.D(_03500_),
    .Q(\cpuregs[15][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _43231_ (.D(_03501_),
    .Q(\cpuregs[15][30] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 _43232_ (.D(_03502_),
    .Q(\cpuregs[15][31] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_4 _43233_ (.D(_03503_),
    .Q(\latched_rd[4] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 _43234_ (.D(_03504_),
    .Q(\cpuregs[7][0] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_1 _43235_ (.D(_03505_),
    .Q(\cpuregs[7][1] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 _43236_ (.D(_03506_),
    .Q(\cpuregs[7][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _43237_ (.D(_03507_),
    .Q(\cpuregs[7][3] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _43238_ (.D(_03508_),
    .Q(\cpuregs[7][4] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 _43239_ (.D(_03509_),
    .Q(\cpuregs[7][5] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _43240_ (.D(_03510_),
    .Q(\cpuregs[7][6] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43241_ (.D(_03511_),
    .Q(\cpuregs[7][7] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _43242_ (.D(_03512_),
    .Q(\cpuregs[7][8] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43243_ (.D(_03513_),
    .Q(\cpuregs[7][9] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43244_ (.D(_03514_),
    .Q(\cpuregs[7][10] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _43245_ (.D(_03515_),
    .Q(\cpuregs[7][11] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 _43246_ (.D(_03516_),
    .Q(\cpuregs[7][12] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43247_ (.D(_03517_),
    .Q(\cpuregs[7][13] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43248_ (.D(_03518_),
    .Q(\cpuregs[7][14] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43249_ (.D(_03519_),
    .Q(\cpuregs[7][15] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _43250_ (.D(_03520_),
    .Q(\cpuregs[7][16] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43251_ (.D(_03521_),
    .Q(\cpuregs[7][17] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43252_ (.D(_03522_),
    .Q(\cpuregs[7][18] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43253_ (.D(_03523_),
    .Q(\cpuregs[7][19] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43254_ (.D(_03524_),
    .Q(\cpuregs[7][20] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _43255_ (.D(_03525_),
    .Q(\cpuregs[7][21] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _43256_ (.D(_03526_),
    .Q(\cpuregs[7][22] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _43257_ (.D(_03527_),
    .Q(\cpuregs[7][23] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _43258_ (.D(_03528_),
    .Q(\cpuregs[7][24] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _43259_ (.D(_03529_),
    .Q(\cpuregs[7][25] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _43260_ (.D(_03530_),
    .Q(\cpuregs[7][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43261_ (.D(_03531_),
    .Q(\cpuregs[7][27] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43262_ (.D(_03532_),
    .Q(\cpuregs[7][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43263_ (.D(_03533_),
    .Q(\cpuregs[7][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _43264_ (.D(_03534_),
    .Q(\cpuregs[7][30] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43265_ (.D(_03535_),
    .Q(\cpuregs[7][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_4 _43266_ (.D(_03536_),
    .Q(net238),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_4 _43267_ (.D(_03537_),
    .Q(net249),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 _43268_ (.D(_03538_),
    .Q(net260),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_4 _43269_ (.D(_03539_),
    .Q(net263),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 _43270_ (.D(_03540_),
    .Q(net264),
    .CLK(clknet_5_15_0_clk));
 sky130_fd_sc_hd__dfxtp_4 _43271_ (.D(_03541_),
    .Q(net265),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_2 _43272_ (.D(_03542_),
    .Q(net266),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _43273_ (.D(_03543_),
    .Q(net267),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__dfxtp_1 _43274_ (.D(_03544_),
    .Q(net268),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__dfxtp_1 _43275_ (.D(_03545_),
    .Q(net269),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_2 _43276_ (.D(_03546_),
    .Q(net239),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_2 _43277_ (.D(_03547_),
    .Q(net240),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_2 _43278_ (.D(_03548_),
    .Q(net241),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 _43279_ (.D(_03549_),
    .Q(net242),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__dfxtp_1 _43280_ (.D(_03550_),
    .Q(net243),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_2 _43281_ (.D(_03551_),
    .Q(net244),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _43282_ (.D(_03552_),
    .Q(net245),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_2 _43283_ (.D(_03553_),
    .Q(net246),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _43284_ (.D(_03554_),
    .Q(net247),
    .CLK(clknet_5_6_0_clk));
 sky130_fd_sc_hd__dfxtp_2 _43285_ (.D(_03555_),
    .Q(net248),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_4 _43286_ (.D(_03556_),
    .Q(net250),
    .CLK(clknet_opt_3_clk));
 sky130_fd_sc_hd__dfxtp_2 _43287_ (.D(_03557_),
    .Q(net251),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 _43288_ (.D(_03558_),
    .Q(net252),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__dfxtp_1 _43289_ (.D(_03559_),
    .Q(net253),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_1 _43290_ (.D(_03560_),
    .Q(net254),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_1 _43291_ (.D(_03561_),
    .Q(net255),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__dfxtp_2 _43292_ (.D(_03562_),
    .Q(net256),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_4 _43293_ (.D(_03563_),
    .Q(net257),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__dfxtp_4 _43294_ (.D(_03564_),
    .Q(net258),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__dfxtp_4 _43295_ (.D(_03565_),
    .Q(net259),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_2 _43296_ (.D(_03566_),
    .Q(net261),
    .CLK(clknet_opt_15_clk));
 sky130_fd_sc_hd__dfxtp_2 _43297_ (.D(_03567_),
    .Q(net262),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__dfxtp_1 _43298_ (.D(_03568_),
    .Q(\cpuregs[19][0] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_1 _43299_ (.D(_03569_),
    .Q(\cpuregs[19][1] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _43300_ (.D(_03570_),
    .Q(\cpuregs[19][2] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 _43301_ (.D(_03571_),
    .Q(\cpuregs[19][3] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43302_ (.D(_03572_),
    .Q(\cpuregs[19][4] ),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__dfxtp_1 _43303_ (.D(_03573_),
    .Q(\cpuregs[19][5] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 _43304_ (.D(_03574_),
    .Q(\cpuregs[19][6] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43305_ (.D(_03575_),
    .Q(\cpuregs[19][7] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _43306_ (.D(_03576_),
    .Q(\cpuregs[19][8] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 _43307_ (.D(_03577_),
    .Q(\cpuregs[19][9] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43308_ (.D(_03578_),
    .Q(\cpuregs[19][10] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 _43309_ (.D(_03579_),
    .Q(\cpuregs[19][11] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 _43310_ (.D(_03580_),
    .Q(\cpuregs[19][12] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43311_ (.D(_03581_),
    .Q(\cpuregs[19][13] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43312_ (.D(_03582_),
    .Q(\cpuregs[19][14] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43313_ (.D(_03583_),
    .Q(\cpuregs[19][15] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43314_ (.D(_03584_),
    .Q(\cpuregs[19][16] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _43315_ (.D(_03585_),
    .Q(\cpuregs[19][17] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43316_ (.D(_03586_),
    .Q(\cpuregs[19][18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _43317_ (.D(_03587_),
    .Q(\cpuregs[19][19] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 _43318_ (.D(_03588_),
    .Q(\cpuregs[19][20] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _43319_ (.D(_03589_),
    .Q(\cpuregs[19][21] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_1 _43320_ (.D(_03590_),
    .Q(\cpuregs[19][22] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_1 _43321_ (.D(_03591_),
    .Q(\cpuregs[19][23] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfxtp_1 _43322_ (.D(_03592_),
    .Q(\cpuregs[19][24] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _43323_ (.D(_03593_),
    .Q(\cpuregs[19][25] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _43324_ (.D(_03594_),
    .Q(\cpuregs[19][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43325_ (.D(_03595_),
    .Q(\cpuregs[19][27] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43326_ (.D(_03596_),
    .Q(\cpuregs[19][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43327_ (.D(_03597_),
    .Q(\cpuregs[19][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _43328_ (.D(_03598_),
    .Q(\cpuregs[19][30] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 _43329_ (.D(_03599_),
    .Q(\cpuregs[19][31] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43330_ (.D(_03600_),
    .Q(\cpuregs[4][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _43331_ (.D(_03601_),
    .Q(\cpuregs[4][1] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _43332_ (.D(_03602_),
    .Q(\cpuregs[4][2] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _43333_ (.D(_03603_),
    .Q(\cpuregs[4][3] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 _43334_ (.D(_03604_),
    .Q(\cpuregs[4][4] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__dfxtp_1 _43335_ (.D(_03605_),
    .Q(\cpuregs[4][5] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _43336_ (.D(_03606_),
    .Q(\cpuregs[4][6] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43337_ (.D(_03607_),
    .Q(\cpuregs[4][7] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _43338_ (.D(_03608_),
    .Q(\cpuregs[4][8] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43339_ (.D(_03609_),
    .Q(\cpuregs[4][9] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43340_ (.D(_03610_),
    .Q(\cpuregs[4][10] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43341_ (.D(_03611_),
    .Q(\cpuregs[4][11] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 _43342_ (.D(_03612_),
    .Q(\cpuregs[4][12] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43343_ (.D(_03613_),
    .Q(\cpuregs[4][13] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 _43344_ (.D(_03614_),
    .Q(\cpuregs[4][14] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 _43345_ (.D(_03615_),
    .Q(\cpuregs[4][15] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 _43346_ (.D(_03616_),
    .Q(\cpuregs[4][16] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43347_ (.D(_03617_),
    .Q(\cpuregs[4][17] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 _43348_ (.D(_03618_),
    .Q(\cpuregs[4][18] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43349_ (.D(_03619_),
    .Q(\cpuregs[4][19] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43350_ (.D(_03620_),
    .Q(\cpuregs[4][20] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _43351_ (.D(_03621_),
    .Q(\cpuregs[4][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__dfxtp_1 _43352_ (.D(_03622_),
    .Q(\cpuregs[4][22] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_1 _43353_ (.D(_03623_),
    .Q(\cpuregs[4][23] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _43354_ (.D(_03624_),
    .Q(\cpuregs[4][24] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _43355_ (.D(_03625_),
    .Q(\cpuregs[4][25] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _43356_ (.D(_03626_),
    .Q(\cpuregs[4][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _43357_ (.D(_03627_),
    .Q(\cpuregs[4][27] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43358_ (.D(_03628_),
    .Q(\cpuregs[4][28] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 _43359_ (.D(_03629_),
    .Q(\cpuregs[4][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfxtp_1 _43360_ (.D(_03630_),
    .Q(\cpuregs[4][30] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43361_ (.D(_03631_),
    .Q(\cpuregs[4][31] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_4 _43362_ (.D(_03632_),
    .Q(net200),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_4 _43363_ (.D(_03633_),
    .Q(net211),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_4 _43364_ (.D(_03634_),
    .Q(net222),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_4 _43365_ (.D(_03635_),
    .Q(net225),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_4 _43366_ (.D(_03636_),
    .Q(net226),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_4 _43367_ (.D(_03637_),
    .Q(net227),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_4 _43368_ (.D(_03638_),
    .Q(net228),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_4 _43369_ (.D(_03639_),
    .Q(net229),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_4 _43370_ (.D(_03640_),
    .Q(net368),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_4 _43371_ (.D(_03641_),
    .Q(net369),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_4 _43372_ (.D(_03642_),
    .Q(net339),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_4 _43373_ (.D(_03643_),
    .Q(net340),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_4 _43374_ (.D(_03644_),
    .Q(net341),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_4 _43375_ (.D(_03645_),
    .Q(net342),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_4 _43376_ (.D(_03646_),
    .Q(net343),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__dfxtp_4 _43377_ (.D(_03647_),
    .Q(net344),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_4 _43378_ (.D(_03648_),
    .Q(net345),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_4 _43379_ (.D(_03649_),
    .Q(net346),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_4 _43380_ (.D(_03650_),
    .Q(net347),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_4 _43381_ (.D(_03651_),
    .Q(net348),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_4 _43382_ (.D(_03652_),
    .Q(net350),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_4 _43383_ (.D(_03653_),
    .Q(net351),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_4 _43384_ (.D(_03654_),
    .Q(net352),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_4 _43385_ (.D(_03655_),
    .Q(net353),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__dfxtp_4 _43386_ (.D(_03656_),
    .Q(net354),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_4 _43387_ (.D(_03657_),
    .Q(net355),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_4 _43388_ (.D(_03658_),
    .Q(net356),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_4 _43389_ (.D(_03659_),
    .Q(net357),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_4 _43390_ (.D(_03660_),
    .Q(net358),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _43391_ (.D(_03661_),
    .Q(net359),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_4 _43392_ (.D(_03662_),
    .Q(net361),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_4 _43393_ (.D(_03663_),
    .Q(net362),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 _43394_ (.D(_03664_),
    .Q(\cpuregs[9][0] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__dfxtp_1 _43395_ (.D(_03665_),
    .Q(\cpuregs[9][1] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 _43396_ (.D(_03666_),
    .Q(\cpuregs[9][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _43397_ (.D(_03667_),
    .Q(\cpuregs[9][3] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 _43398_ (.D(_03668_),
    .Q(\cpuregs[9][4] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__dfxtp_1 _43399_ (.D(_03669_),
    .Q(\cpuregs[9][5] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _43400_ (.D(_03670_),
    .Q(\cpuregs[9][6] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43401_ (.D(_03671_),
    .Q(\cpuregs[9][7] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__dfxtp_1 _43402_ (.D(_03672_),
    .Q(\cpuregs[9][8] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 _43403_ (.D(_03673_),
    .Q(\cpuregs[9][9] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43404_ (.D(_03674_),
    .Q(\cpuregs[9][10] ),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__dfxtp_1 _43405_ (.D(_03675_),
    .Q(\cpuregs[9][11] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 _43406_ (.D(_03676_),
    .Q(\cpuregs[9][12] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 _43407_ (.D(_03677_),
    .Q(\cpuregs[9][13] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43408_ (.D(_03678_),
    .Q(\cpuregs[9][14] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43409_ (.D(_03679_),
    .Q(\cpuregs[9][15] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43410_ (.D(_03680_),
    .Q(\cpuregs[9][16] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _43411_ (.D(_03681_),
    .Q(\cpuregs[9][17] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43412_ (.D(_03682_),
    .Q(\cpuregs[9][18] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 _43413_ (.D(_03683_),
    .Q(\cpuregs[9][19] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _43414_ (.D(_03684_),
    .Q(\cpuregs[9][20] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43415_ (.D(_03685_),
    .Q(\cpuregs[9][21] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 _43416_ (.D(_03686_),
    .Q(\cpuregs[9][22] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 _43417_ (.D(_03687_),
    .Q(\cpuregs[9][23] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__dfxtp_1 _43418_ (.D(_03688_),
    .Q(\cpuregs[9][24] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43419_ (.D(_03689_),
    .Q(\cpuregs[9][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__dfxtp_1 _43420_ (.D(_03690_),
    .Q(\cpuregs[9][26] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43421_ (.D(_03691_),
    .Q(\cpuregs[9][27] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43422_ (.D(_03692_),
    .Q(\cpuregs[9][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43423_ (.D(_03693_),
    .Q(\cpuregs[9][29] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43424_ (.D(_03694_),
    .Q(\cpuregs[9][30] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 _43425_ (.D(_03695_),
    .Q(\cpuregs[9][31] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 _43426_ (.D(_03696_),
    .Q(\cpuregs[6][0] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_1 _43427_ (.D(_03697_),
    .Q(\cpuregs[6][1] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 _43428_ (.D(_03698_),
    .Q(\cpuregs[6][2] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__dfxtp_1 _43429_ (.D(_03699_),
    .Q(\cpuregs[6][3] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__dfxtp_1 _43430_ (.D(_03700_),
    .Q(\cpuregs[6][4] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__dfxtp_1 _43431_ (.D(_03701_),
    .Q(\cpuregs[6][5] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__dfxtp_1 _43432_ (.D(_03702_),
    .Q(\cpuregs[6][6] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43433_ (.D(_03703_),
    .Q(\cpuregs[6][7] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 _43434_ (.D(_03704_),
    .Q(\cpuregs[6][8] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 _43435_ (.D(_03705_),
    .Q(\cpuregs[6][9] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43436_ (.D(_03706_),
    .Q(\cpuregs[6][10] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 _43437_ (.D(_03707_),
    .Q(\cpuregs[6][11] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 _43438_ (.D(_03708_),
    .Q(\cpuregs[6][12] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 _43439_ (.D(_03709_),
    .Q(\cpuregs[6][13] ),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__dfxtp_1 _43440_ (.D(_03710_),
    .Q(\cpuregs[6][14] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43441_ (.D(_03711_),
    .Q(\cpuregs[6][15] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 _43442_ (.D(_03712_),
    .Q(\cpuregs[6][16] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 _43443_ (.D(_03713_),
    .Q(\cpuregs[6][17] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 _43444_ (.D(_03714_),
    .Q(\cpuregs[6][18] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 _43445_ (.D(_03715_),
    .Q(\cpuregs[6][19] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 _43446_ (.D(_03716_),
    .Q(\cpuregs[6][20] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _43447_ (.D(_03717_),
    .Q(\cpuregs[6][21] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_1 _43448_ (.D(_03718_),
    .Q(\cpuregs[6][22] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__dfxtp_1 _43449_ (.D(_03719_),
    .Q(\cpuregs[6][23] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__dfxtp_1 _43450_ (.D(_03720_),
    .Q(\cpuregs[6][24] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _43451_ (.D(_03721_),
    .Q(\cpuregs[6][25] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfxtp_1 _43452_ (.D(_03722_),
    .Q(\cpuregs[6][26] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 _43453_ (.D(_03723_),
    .Q(\cpuregs[6][27] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43454_ (.D(_03724_),
    .Q(\cpuregs[6][28] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfxtp_1 _43455_ (.D(_03725_),
    .Q(\cpuregs[6][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 _43456_ (.D(_03726_),
    .Q(\cpuregs[6][30] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43457_ (.D(_03727_),
    .Q(\cpuregs[6][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfxtp_1 _43458_ (.D(_03728_),
    .Q(\pcpi_mul.active[0] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_4 _43459_ (.D(_03729_),
    .Q(\pcpi_mul.active[1] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_4 _43460_ (.D(_03730_),
    .Q(net408),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 _43461_ (.D(_03731_),
    .Q(\count_cycle[0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 _43462_ (.D(_03732_),
    .Q(\count_cycle[1] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 _43463_ (.D(_03733_),
    .Q(\count_cycle[2] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 _43464_ (.D(_03734_),
    .Q(\count_cycle[3] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43465_ (.D(_03735_),
    .Q(\count_cycle[4] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43466_ (.D(_03736_),
    .Q(\count_cycle[5] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43467_ (.D(_03737_),
    .Q(\count_cycle[6] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43468_ (.D(_03738_),
    .Q(\count_cycle[7] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _43469_ (.D(_03739_),
    .Q(\count_cycle[8] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfxtp_1 _43470_ (.D(_03740_),
    .Q(\count_cycle[9] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _43471_ (.D(_03741_),
    .Q(\count_cycle[10] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _43472_ (.D(_03742_),
    .Q(\count_cycle[11] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _43473_ (.D(_03743_),
    .Q(\count_cycle[12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43474_ (.D(_03744_),
    .Q(\count_cycle[13] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43475_ (.D(_03745_),
    .Q(\count_cycle[14] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43476_ (.D(_03746_),
    .Q(\count_cycle[15] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43477_ (.D(_03747_),
    .Q(\count_cycle[16] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 _43478_ (.D(_03748_),
    .Q(\count_cycle[17] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43479_ (.D(_03749_),
    .Q(\count_cycle[18] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43480_ (.D(_03750_),
    .Q(\count_cycle[19] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43481_ (.D(_03751_),
    .Q(\count_cycle[20] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43482_ (.D(_03752_),
    .Q(\count_cycle[21] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43483_ (.D(_03753_),
    .Q(\count_cycle[22] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43484_ (.D(_03754_),
    .Q(\count_cycle[23] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43485_ (.D(_03755_),
    .Q(\count_cycle[24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43486_ (.D(_03756_),
    .Q(\count_cycle[25] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43487_ (.D(_03757_),
    .Q(\count_cycle[26] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43488_ (.D(_03758_),
    .Q(\count_cycle[27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43489_ (.D(_03759_),
    .Q(\count_cycle[28] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _43490_ (.D(_03760_),
    .Q(\count_cycle[29] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 _43491_ (.D(_03761_),
    .Q(\count_cycle[30] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 _43492_ (.D(_03762_),
    .Q(\count_cycle[31] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 _43493_ (.D(_03763_),
    .Q(\count_cycle[32] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 _43494_ (.D(_03764_),
    .Q(\count_cycle[33] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 _43495_ (.D(_03765_),
    .Q(\count_cycle[34] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 _43496_ (.D(_03766_),
    .Q(\count_cycle[35] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _43497_ (.D(_03767_),
    .Q(\count_cycle[36] ),
    .CLK(clknet_5_25_0_clk));
 sky130_fd_sc_hd__dfxtp_1 _43498_ (.D(_03768_),
    .Q(\count_cycle[37] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43499_ (.D(_03769_),
    .Q(\count_cycle[38] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43500_ (.D(_03770_),
    .Q(\count_cycle[39] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43501_ (.D(_03771_),
    .Q(\count_cycle[40] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43502_ (.D(_03772_),
    .Q(\count_cycle[41] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43503_ (.D(_03773_),
    .Q(\count_cycle[42] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _43504_ (.D(_03774_),
    .Q(\count_cycle[43] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _43505_ (.D(_03775_),
    .Q(\count_cycle[44] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _43506_ (.D(_03776_),
    .Q(\count_cycle[45] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _43507_ (.D(_03777_),
    .Q(\count_cycle[46] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _43508_ (.D(_03778_),
    .Q(\count_cycle[47] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__dfxtp_1 _43509_ (.D(_03779_),
    .Q(\count_cycle[48] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _43510_ (.D(_03780_),
    .Q(\count_cycle[49] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43511_ (.D(_03781_),
    .Q(\count_cycle[50] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43512_ (.D(_03782_),
    .Q(\count_cycle[51] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43513_ (.D(_03783_),
    .Q(\count_cycle[52] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43514_ (.D(_03784_),
    .Q(\count_cycle[53] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43515_ (.D(_03785_),
    .Q(\count_cycle[54] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43516_ (.D(_03786_),
    .Q(\count_cycle[55] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43517_ (.D(_03787_),
    .Q(\count_cycle[56] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43518_ (.D(_03788_),
    .Q(\count_cycle[57] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43519_ (.D(_03789_),
    .Q(\count_cycle[58] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43520_ (.D(_03790_),
    .Q(\count_cycle[59] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43521_ (.D(_03791_),
    .Q(\count_cycle[60] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43522_ (.D(_03792_),
    .Q(\count_cycle[61] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 _43523_ (.D(_03793_),
    .Q(\count_cycle[62] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 _43524_ (.D(_03794_),
    .Q(\count_cycle[63] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43525_ (.D(_03795_),
    .Q(\timer[0] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 _43526_ (.D(_03796_),
    .Q(\timer[1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _43527_ (.D(_03797_),
    .Q(\timer[2] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _43528_ (.D(_03798_),
    .Q(\timer[3] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 _43529_ (.D(_03799_),
    .Q(\timer[4] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 _43530_ (.D(_03800_),
    .Q(\timer[5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 _43531_ (.D(_03801_),
    .Q(\timer[6] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 _43532_ (.D(_03802_),
    .Q(\timer[7] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 _43533_ (.D(_03803_),
    .Q(\timer[8] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 _43534_ (.D(_03804_),
    .Q(\timer[9] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _43535_ (.D(_03805_),
    .Q(\timer[10] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 _43536_ (.D(_03806_),
    .Q(\timer[11] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _43537_ (.D(_03807_),
    .Q(\timer[12] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _43538_ (.D(_03808_),
    .Q(\timer[13] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _43539_ (.D(_03809_),
    .Q(\timer[14] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43540_ (.D(_03810_),
    .Q(\timer[15] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _43541_ (.D(_03811_),
    .Q(\timer[16] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _43542_ (.D(_03812_),
    .Q(\timer[17] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 _43543_ (.D(_03813_),
    .Q(\timer[18] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 _43544_ (.D(_03814_),
    .Q(\timer[19] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _43545_ (.D(_03815_),
    .Q(\timer[20] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _43546_ (.D(_03816_),
    .Q(\timer[21] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _43547_ (.D(_03817_),
    .Q(\timer[22] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43548_ (.D(_03818_),
    .Q(\timer[23] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43549_ (.D(_03819_),
    .Q(\timer[24] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43550_ (.D(_03820_),
    .Q(\timer[25] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 _43551_ (.D(_03821_),
    .Q(\timer[26] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 _43552_ (.D(_03822_),
    .Q(\timer[27] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43553_ (.D(_03823_),
    .Q(\timer[28] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 _43554_ (.D(_03824_),
    .Q(\timer[29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 _43555_ (.D(_03825_),
    .Q(\timer[30] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 _43556_ (.D(_03826_),
    .Q(\timer[31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_2 _43557_ (.D(_03827_),
    .Q(pcpi_timeout),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43558_ (.D(_03828_),
    .Q(decoder_pseudo_trigger),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_4 _43559_ (.D(_03829_),
    .Q(is_compare),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 _43560_ (.D(_03830_),
    .Q(do_waitirq),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_4 _43561_ (.D(_03831_),
    .Q(net237),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_4 _43562_ (.D(_03832_),
    .Q(net370),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_4 _43563_ (.D(_03833_),
    .Q(net102),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _43564_ (.D(_03834_),
    .Q(net113),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_4 _43565_ (.D(_03835_),
    .Q(net124),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_4 _43566_ (.D(_03836_),
    .Q(net127),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_4 _43567_ (.D(_03837_),
    .Q(net128),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_4 _43568_ (.D(_03838_),
    .Q(net129),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_4 _43569_ (.D(_03839_),
    .Q(net130),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_2 _43570_ (.D(_03840_),
    .Q(net131),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_4 _43571_ (.D(_03841_),
    .Q(net132),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_4 _43572_ (.D(_03842_),
    .Q(net133),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_4 _43573_ (.D(_03843_),
    .Q(net103),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__dfxtp_4 _43574_ (.D(_03844_),
    .Q(net104),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_4 _43575_ (.D(_03845_),
    .Q(net105),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_4 _43576_ (.D(_03846_),
    .Q(net106),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 _43577_ (.D(_03847_),
    .Q(net107),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _43578_ (.D(_03848_),
    .Q(net108),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_4 _43579_ (.D(_03849_),
    .Q(net109),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_4 _43580_ (.D(_03850_),
    .Q(net110),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__dfxtp_2 _43581_ (.D(_03851_),
    .Q(net111),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_4 _43582_ (.D(_03852_),
    .Q(net112),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_4 _43583_ (.D(_03853_),
    .Q(net114),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_4 _43584_ (.D(_03854_),
    .Q(net115),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_2 _43585_ (.D(_03855_),
    .Q(net116),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__dfxtp_4 _43586_ (.D(_03856_),
    .Q(net117),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_4 _43587_ (.D(_03857_),
    .Q(net118),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _43588_ (.D(_03858_),
    .Q(net119),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__dfxtp_4 _43589_ (.D(_03859_),
    .Q(net120),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_4 _43590_ (.D(_03860_),
    .Q(net121),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_4 _43591_ (.D(_03861_),
    .Q(net122),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_4 _43592_ (.D(_03862_),
    .Q(net123),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_2 _43593_ (.D(_03863_),
    .Q(net125),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_4 _43594_ (.D(_03864_),
    .Q(net126),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 _43595_ (.D(_03865_),
    .Q(\count_instr[0] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 _43596_ (.D(_03866_),
    .Q(\count_instr[1] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 _43597_ (.D(_03867_),
    .Q(\count_instr[2] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfxtp_1 _43598_ (.D(_03868_),
    .Q(\count_instr[3] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 _43599_ (.D(_03869_),
    .Q(\count_instr[4] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 _43600_ (.D(_03870_),
    .Q(\count_instr[5] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43601_ (.D(_03871_),
    .Q(\count_instr[6] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43602_ (.D(_03872_),
    .Q(\count_instr[7] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43603_ (.D(_03873_),
    .Q(\count_instr[8] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__dfxtp_1 _43604_ (.D(_03874_),
    .Q(\count_instr[9] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _43605_ (.D(_03875_),
    .Q(\count_instr[10] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__dfxtp_1 _43606_ (.D(_03876_),
    .Q(\count_instr[11] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43607_ (.D(_03877_),
    .Q(\count_instr[12] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _43608_ (.D(_03878_),
    .Q(\count_instr[13] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43609_ (.D(_03879_),
    .Q(\count_instr[14] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43610_ (.D(_03880_),
    .Q(\count_instr[15] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43611_ (.D(_03881_),
    .Q(\count_instr[16] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43612_ (.D(_03882_),
    .Q(\count_instr[17] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43613_ (.D(_03883_),
    .Q(\count_instr[18] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43614_ (.D(_03884_),
    .Q(\count_instr[19] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43615_ (.D(_03885_),
    .Q(\count_instr[20] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43616_ (.D(_03886_),
    .Q(\count_instr[21] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43617_ (.D(_03887_),
    .Q(\count_instr[22] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43618_ (.D(_03888_),
    .Q(\count_instr[23] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 _43619_ (.D(_03889_),
    .Q(\count_instr[24] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 _43620_ (.D(_03890_),
    .Q(\count_instr[25] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43621_ (.D(_03891_),
    .Q(\count_instr[26] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43622_ (.D(_03892_),
    .Q(\count_instr[27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43623_ (.D(_03893_),
    .Q(\count_instr[28] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43624_ (.D(_03894_),
    .Q(\count_instr[29] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43625_ (.D(_03895_),
    .Q(\count_instr[30] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 _43626_ (.D(_03896_),
    .Q(\count_instr[31] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43627_ (.D(_03897_),
    .Q(\count_instr[32] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43628_ (.D(_03898_),
    .Q(\count_instr[33] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43629_ (.D(_03899_),
    .Q(\count_instr[34] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 _43630_ (.D(_03900_),
    .Q(\count_instr[35] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 _43631_ (.D(_03901_),
    .Q(\count_instr[36] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__dfxtp_1 _43632_ (.D(_03902_),
    .Q(\count_instr[37] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43633_ (.D(_03903_),
    .Q(\count_instr[38] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43634_ (.D(_03904_),
    .Q(\count_instr[39] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43635_ (.D(_03905_),
    .Q(\count_instr[40] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 _43636_ (.D(_03906_),
    .Q(\count_instr[41] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__dfxtp_1 _43637_ (.D(_03907_),
    .Q(\count_instr[42] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _43638_ (.D(_03908_),
    .Q(\count_instr[43] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _43639_ (.D(_03909_),
    .Q(\count_instr[44] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__dfxtp_1 _43640_ (.D(_03910_),
    .Q(\count_instr[45] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43641_ (.D(_03911_),
    .Q(\count_instr[46] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 _43642_ (.D(_03912_),
    .Q(\count_instr[47] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43643_ (.D(_03913_),
    .Q(\count_instr[48] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43644_ (.D(_03914_),
    .Q(\count_instr[49] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43645_ (.D(_03915_),
    .Q(\count_instr[50] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43646_ (.D(_03916_),
    .Q(\count_instr[51] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 _43647_ (.D(_03917_),
    .Q(\count_instr[52] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43648_ (.D(_03918_),
    .Q(\count_instr[53] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43649_ (.D(_03919_),
    .Q(\count_instr[54] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43650_ (.D(_03920_),
    .Q(\count_instr[55] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 _43651_ (.D(_03921_),
    .Q(\count_instr[56] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43652_ (.D(_03922_),
    .Q(\count_instr[57] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43653_ (.D(_03923_),
    .Q(\count_instr[58] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43654_ (.D(_03924_),
    .Q(\count_instr[59] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43655_ (.D(_03925_),
    .Q(\count_instr[60] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 _43656_ (.D(_03926_),
    .Q(\count_instr[61] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 _43657_ (.D(_03927_),
    .Q(\count_instr[62] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 _43658_ (.D(_03928_),
    .Q(\count_instr[63] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_2 _43659_ (.D(_03929_),
    .Q(\reg_pc[1] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_2 _43660_ (.D(_03930_),
    .Q(\reg_pc[2] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 _43661_ (.D(_03931_),
    .Q(\reg_pc[3] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 _43662_ (.D(_03932_),
    .Q(\reg_pc[4] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 _43663_ (.D(_03933_),
    .Q(\reg_pc[5] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 _43664_ (.D(_03934_),
    .Q(\reg_pc[6] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_2 _43665_ (.D(_03935_),
    .Q(\reg_pc[7] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__dfxtp_1 _43666_ (.D(_03936_),
    .Q(\reg_pc[8] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_2 _43667_ (.D(_03937_),
    .Q(\reg_pc[9] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 _43668_ (.D(_03938_),
    .Q(\reg_pc[10] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_2 _43669_ (.D(_03939_),
    .Q(\reg_pc[11] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_1 _43670_ (.D(_03940_),
    .Q(\reg_pc[12] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_2 _43671_ (.D(_03941_),
    .Q(\reg_pc[13] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_2 _43672_ (.D(_03942_),
    .Q(\reg_pc[14] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _43673_ (.D(_03943_),
    .Q(\reg_pc[15] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_1 _43674_ (.D(_03944_),
    .Q(\reg_pc[16] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_2 _43675_ (.D(_03945_),
    .Q(\reg_pc[17] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__dfxtp_4 _43676_ (.D(_03946_),
    .Q(\reg_pc[18] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43677_ (.D(_03947_),
    .Q(\reg_pc[19] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_4 _43678_ (.D(_03948_),
    .Q(\reg_pc[20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_2 _43679_ (.D(_03949_),
    .Q(\reg_pc[21] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_4 _43680_ (.D(_03950_),
    .Q(\reg_pc[22] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_2 _43681_ (.D(_03951_),
    .Q(\reg_pc[23] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _43682_ (.D(_03952_),
    .Q(\reg_pc[24] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _43683_ (.D(_03953_),
    .Q(\reg_pc[25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _43684_ (.D(_03954_),
    .Q(\reg_pc[26] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_4 _43685_ (.D(_03955_),
    .Q(\reg_pc[27] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_4 _43686_ (.D(_03956_),
    .Q(\reg_pc[28] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _43687_ (.D(_03957_),
    .Q(\reg_pc[29] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_4 _43688_ (.D(_03958_),
    .Q(\reg_pc[30] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_2 _43689_ (.D(_03959_),
    .Q(\reg_pc[31] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _43690_ (.D(_03960_),
    .Q(\reg_next_pc[1] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 _43691_ (.D(_03961_),
    .Q(\reg_next_pc[2] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 _43692_ (.D(_03962_),
    .Q(\reg_next_pc[3] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 _43693_ (.D(_03963_),
    .Q(\reg_next_pc[4] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 _43694_ (.D(_03964_),
    .Q(\reg_next_pc[5] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 _43695_ (.D(_03965_),
    .Q(\reg_next_pc[6] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 _43696_ (.D(_03966_),
    .Q(\reg_next_pc[7] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__dfxtp_1 _43697_ (.D(_03967_),
    .Q(\reg_next_pc[8] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__dfxtp_1 _43698_ (.D(_03968_),
    .Q(\reg_next_pc[9] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__dfxtp_1 _43699_ (.D(_03969_),
    .Q(\reg_next_pc[10] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_1 _43700_ (.D(_03970_),
    .Q(\reg_next_pc[11] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_1 _43701_ (.D(_03971_),
    .Q(\reg_next_pc[12] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_2 _43702_ (.D(_03972_),
    .Q(\reg_next_pc[13] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43703_ (.D(_03973_),
    .Q(\reg_next_pc[14] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43704_ (.D(_03974_),
    .Q(\reg_next_pc[15] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _43705_ (.D(_03975_),
    .Q(\reg_next_pc[16] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _43706_ (.D(_03976_),
    .Q(\reg_next_pc[17] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 _43707_ (.D(_03977_),
    .Q(\reg_next_pc[18] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _43708_ (.D(_03978_),
    .Q(\reg_next_pc[19] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _43709_ (.D(_03979_),
    .Q(\reg_next_pc[20] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__dfxtp_1 _43710_ (.D(_03980_),
    .Q(\reg_next_pc[21] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43711_ (.D(_03981_),
    .Q(\reg_next_pc[22] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__dfxtp_1 _43712_ (.D(_03982_),
    .Q(\reg_next_pc[23] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_1 _43713_ (.D(_03983_),
    .Q(\reg_next_pc[24] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _43714_ (.D(_03984_),
    .Q(\reg_next_pc[25] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _43715_ (.D(_03985_),
    .Q(\reg_next_pc[26] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _43716_ (.D(_03986_),
    .Q(\reg_next_pc[27] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _43717_ (.D(_03987_),
    .Q(\reg_next_pc[28] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__dfxtp_2 _43718_ (.D(_03988_),
    .Q(\reg_next_pc[29] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__dfxtp_2 _43719_ (.D(_03989_),
    .Q(\reg_next_pc[30] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__dfxtp_1 _43720_ (.D(_03990_),
    .Q(\reg_next_pc[31] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__dfxtp_2 _43721_ (.D(_03991_),
    .Q(mem_do_rdata),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 _43722_ (.D(_03992_),
    .Q(mem_do_wdata),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 _43723_ (.D(_03993_),
    .Q(\pcpi_timeout_counter[0] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43724_ (.D(_03994_),
    .Q(\pcpi_timeout_counter[1] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43725_ (.D(_03995_),
    .Q(\pcpi_timeout_counter[2] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _43726_ (.D(_03996_),
    .Q(\pcpi_timeout_counter[3] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_1 _43727_ (.D(_03997_),
    .Q(instr_beq),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _43728_ (.D(_03998_),
    .Q(instr_bne),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _43729_ (.D(_03999_),
    .Q(instr_blt),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _43730_ (.D(_04000_),
    .Q(instr_bge),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 _43731_ (.D(_04001_),
    .Q(instr_bltu),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _43732_ (.D(_04002_),
    .Q(instr_bgeu),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43733_ (.D(_04003_),
    .Q(instr_addi),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _43734_ (.D(_04004_),
    .Q(instr_slti),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 _43735_ (.D(_04005_),
    .Q(instr_sltiu),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_2 _43736_ (.D(_04006_),
    .Q(instr_xori),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_2 _43737_ (.D(_04007_),
    .Q(instr_ori),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _43738_ (.D(_04008_),
    .Q(instr_andi),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43739_ (.D(_04009_),
    .Q(instr_add),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_4 _43740_ (.D(_04010_),
    .Q(instr_sub),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 _43741_ (.D(_04011_),
    .Q(instr_sll),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _43742_ (.D(_04012_),
    .Q(instr_slt),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _43743_ (.D(_04013_),
    .Q(instr_sltu),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_2 _43744_ (.D(_04014_),
    .Q(instr_xor),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 _43745_ (.D(_04015_),
    .Q(instr_srl),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 _43746_ (.D(_04016_),
    .Q(instr_sra),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_2 _43747_ (.D(_04017_),
    .Q(instr_or),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfxtp_2 _43748_ (.D(_04018_),
    .Q(instr_and),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfxtp_1 _43749_ (.D(_04019_),
    .Q(\decoded_rs1[0] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 _43750_ (.D(_04020_),
    .Q(\decoded_rs1[1] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 _43751_ (.D(_04021_),
    .Q(\decoded_rs1[2] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 _43752_ (.D(_04022_),
    .Q(\decoded_rs1[3] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_4 _43753_ (.D(_04023_),
    .Q(is_beq_bne_blt_bge_bltu_bgeu),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 _43754_ (.D(_04024_),
    .Q(net166),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 _43755_ (.D(_04025_),
    .Q(\irq_mask[0] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 _43756_ (.D(_04026_),
    .Q(\irq_mask[1] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _43757_ (.D(_04027_),
    .Q(\irq_mask[2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _43758_ (.D(_04028_),
    .Q(\irq_mask[3] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _43759_ (.D(_04029_),
    .Q(\irq_mask[4] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _43760_ (.D(_04030_),
    .Q(\irq_mask[5] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43761_ (.D(_04031_),
    .Q(\irq_mask[6] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _43762_ (.D(_04032_),
    .Q(\irq_mask[7] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43763_ (.D(_04033_),
    .Q(\irq_mask[8] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_2 _43764_ (.D(_04034_),
    .Q(\irq_mask[9] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 _43765_ (.D(_04035_),
    .Q(\irq_mask[10] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_1 _43766_ (.D(_04036_),
    .Q(\irq_mask[11] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_1 _43767_ (.D(_04037_),
    .Q(\irq_mask[12] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _43768_ (.D(_04038_),
    .Q(\irq_mask[13] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 _43769_ (.D(_04039_),
    .Q(\irq_mask[14] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _43770_ (.D(_04040_),
    .Q(\irq_mask[15] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_2 _43771_ (.D(_04041_),
    .Q(\irq_mask[16] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _43772_ (.D(_04042_),
    .Q(\irq_mask[17] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 _43773_ (.D(_04043_),
    .Q(\irq_mask[18] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _43774_ (.D(_04044_),
    .Q(\irq_mask[19] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 _43775_ (.D(_04045_),
    .Q(\irq_mask[20] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__dfxtp_1 _43776_ (.D(_04046_),
    .Q(\irq_mask[21] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _43777_ (.D(_04047_),
    .Q(\irq_mask[22] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_2 _43778_ (.D(_04048_),
    .Q(\irq_mask[23] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43779_ (.D(_04049_),
    .Q(\irq_mask[24] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_2 _43780_ (.D(_04050_),
    .Q(\irq_mask[25] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 _43781_ (.D(_04051_),
    .Q(\irq_mask[26] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43782_ (.D(_04052_),
    .Q(\irq_mask[27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43783_ (.D(_04053_),
    .Q(\irq_mask[28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 _43784_ (.D(_04054_),
    .Q(\irq_mask[29] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _43785_ (.D(_04055_),
    .Q(\irq_mask[30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 _43786_ (.D(_04056_),
    .Q(\irq_mask[31] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 _43787_ (.D(_04057_),
    .Q(mem_do_prefetch),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 _43788_ (.D(_04058_),
    .Q(mem_do_rinst),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 _43789_ (.D(_04059_),
    .Q(\irq_state[0] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_4 _43790_ (.D(_04060_),
    .Q(\irq_state[1] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_4 _43791_ (.D(_04061_),
    .Q(latched_store),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_4 _43792_ (.D(_04062_),
    .Q(latched_stalu),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_4 _43793_ (.D(_04063_),
    .Q(\pcpi_mul.rs2[32] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_2 _43794_ (.D(_04064_),
    .Q(\pcpi_mul.rs1[32] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 _43795_ (.D(_04065_),
    .Q(irq_delay),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 _43796_ (.D(_04066_),
    .Q(\decoded_rs1[4] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_2 _43797_ (.D(_04067_),
    .Q(\mem_state[0] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_2 _43798_ (.D(_04068_),
    .Q(\mem_state[1] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_4 _43799_ (.D(_04069_),
    .Q(latched_branch),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_2 _43800_ (.D(_04070_),
    .Q(latched_is_lh),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_2 _43801_ (.D(_04071_),
    .Q(latched_is_lb),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 _43802_ (.D(_04072_),
    .Q(irq_active),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8828 ();
 sky130_fd_sc_hd__clkbuf_8 input1 (.A(irq[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(irq[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(irq[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input4 (.A(irq[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_8 input5 (.A(irq[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input6 (.A(irq[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(irq[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(irq[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(irq[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(irq[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(irq[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(irq[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(irq[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(irq[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(irq[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(irq[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(irq[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input18 (.A(irq[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(irq[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(irq[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(irq[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_6 input22 (.A(irq[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_6 input23 (.A(irq[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_6 input24 (.A(irq[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(irq[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(irq[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(irq[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(irq[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_6 input29 (.A(irq[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(irq[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(irq[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(irq[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_6 input33 (.A(mem_rdata[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(mem_rdata[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_6 input35 (.A(mem_rdata[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(mem_rdata[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input37 (.A(mem_rdata[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_6 input38 (.A(mem_rdata[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(mem_rdata[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_6 input40 (.A(mem_rdata[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_6 input41 (.A(mem_rdata[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_6 input42 (.A(mem_rdata[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(mem_rdata[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_8 input44 (.A(mem_rdata[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(mem_rdata[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(mem_rdata[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_8 input47 (.A(mem_rdata[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(mem_rdata[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_6 input49 (.A(mem_rdata[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 input50 (.A(mem_rdata[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_6 input51 (.A(mem_rdata[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_6 input52 (.A(mem_rdata[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_4 input53 (.A(mem_rdata[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_6 input54 (.A(mem_rdata[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_6 input55 (.A(mem_rdata[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(mem_rdata[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_6 input57 (.A(mem_rdata[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_6 input58 (.A(mem_rdata[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_8 input59 (.A(mem_rdata[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(mem_rdata[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(mem_rdata[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_6 input62 (.A(mem_rdata[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_8 input63 (.A(mem_rdata[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(mem_rdata[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(mem_ready),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(pcpi_rd[0]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(pcpi_rd[10]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(pcpi_rd[11]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(pcpi_rd[12]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(pcpi_rd[13]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(pcpi_rd[14]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(pcpi_rd[15]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(pcpi_rd[16]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(pcpi_rd[17]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(pcpi_rd[18]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(pcpi_rd[19]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(pcpi_rd[1]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(pcpi_rd[20]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(pcpi_rd[21]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(pcpi_rd[22]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(pcpi_rd[23]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(pcpi_rd[24]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(pcpi_rd[25]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(pcpi_rd[26]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(pcpi_rd[27]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(pcpi_rd[28]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(pcpi_rd[29]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(pcpi_rd[2]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(pcpi_rd[30]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(pcpi_rd[31]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(pcpi_rd[3]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(pcpi_rd[4]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(pcpi_rd[5]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(pcpi_rd[6]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(pcpi_rd[7]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(pcpi_rd[8]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(pcpi_rd[9]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(pcpi_ready),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(pcpi_wait),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(pcpi_wr),
    .X(net100));
 sky130_fd_sc_hd__buf_4 input101 (.A(resetn),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(eoi[0]));
 sky130_fd_sc_hd__clkbuf_2 output103 (.A(net103),
    .X(eoi[10]));
 sky130_fd_sc_hd__clkbuf_2 output104 (.A(net104),
    .X(eoi[11]));
 sky130_fd_sc_hd__clkbuf_2 output105 (.A(net105),
    .X(eoi[12]));
 sky130_fd_sc_hd__clkbuf_2 output106 (.A(net106),
    .X(eoi[13]));
 sky130_fd_sc_hd__clkbuf_2 output107 (.A(net107),
    .X(eoi[14]));
 sky130_fd_sc_hd__clkbuf_2 output108 (.A(net108),
    .X(eoi[15]));
 sky130_fd_sc_hd__clkbuf_2 output109 (.A(net109),
    .X(eoi[16]));
 sky130_fd_sc_hd__clkbuf_2 output110 (.A(net110),
    .X(eoi[17]));
 sky130_fd_sc_hd__clkbuf_2 output111 (.A(net111),
    .X(eoi[18]));
 sky130_fd_sc_hd__clkbuf_2 output112 (.A(net112),
    .X(eoi[19]));
 sky130_fd_sc_hd__clkbuf_2 output113 (.A(net113),
    .X(eoi[1]));
 sky130_fd_sc_hd__clkbuf_2 output114 (.A(net114),
    .X(eoi[20]));
 sky130_fd_sc_hd__clkbuf_2 output115 (.A(net115),
    .X(eoi[21]));
 sky130_fd_sc_hd__clkbuf_2 output116 (.A(net116),
    .X(eoi[22]));
 sky130_fd_sc_hd__clkbuf_2 output117 (.A(net117),
    .X(eoi[23]));
 sky130_fd_sc_hd__clkbuf_2 output118 (.A(net118),
    .X(eoi[24]));
 sky130_fd_sc_hd__clkbuf_2 output119 (.A(net119),
    .X(eoi[25]));
 sky130_fd_sc_hd__clkbuf_2 output120 (.A(net120),
    .X(eoi[26]));
 sky130_fd_sc_hd__clkbuf_2 output121 (.A(net121),
    .X(eoi[27]));
 sky130_fd_sc_hd__clkbuf_2 output122 (.A(net122),
    .X(eoi[28]));
 sky130_fd_sc_hd__clkbuf_2 output123 (.A(net123),
    .X(eoi[29]));
 sky130_fd_sc_hd__clkbuf_2 output124 (.A(net124),
    .X(eoi[2]));
 sky130_fd_sc_hd__clkbuf_2 output125 (.A(net125),
    .X(eoi[30]));
 sky130_fd_sc_hd__clkbuf_2 output126 (.A(net126),
    .X(eoi[31]));
 sky130_fd_sc_hd__clkbuf_2 output127 (.A(net127),
    .X(eoi[3]));
 sky130_fd_sc_hd__clkbuf_2 output128 (.A(net128),
    .X(eoi[4]));
 sky130_fd_sc_hd__clkbuf_2 output129 (.A(net129),
    .X(eoi[5]));
 sky130_fd_sc_hd__clkbuf_2 output130 (.A(net130),
    .X(eoi[6]));
 sky130_fd_sc_hd__clkbuf_2 output131 (.A(net131),
    .X(eoi[7]));
 sky130_fd_sc_hd__clkbuf_2 output132 (.A(net132),
    .X(eoi[8]));
 sky130_fd_sc_hd__clkbuf_2 output133 (.A(net133),
    .X(eoi[9]));
 sky130_fd_sc_hd__clkbuf_2 output134 (.A(net134),
    .X(mem_addr[0]));
 sky130_fd_sc_hd__clkbuf_2 output135 (.A(net135),
    .X(mem_addr[10]));
 sky130_fd_sc_hd__clkbuf_2 output136 (.A(net136),
    .X(mem_addr[11]));
 sky130_fd_sc_hd__clkbuf_2 output137 (.A(net137),
    .X(mem_addr[12]));
 sky130_fd_sc_hd__clkbuf_2 output138 (.A(net138),
    .X(mem_addr[13]));
 sky130_fd_sc_hd__clkbuf_2 output139 (.A(net139),
    .X(mem_addr[14]));
 sky130_fd_sc_hd__clkbuf_2 output140 (.A(net140),
    .X(mem_addr[15]));
 sky130_fd_sc_hd__clkbuf_2 output141 (.A(net141),
    .X(mem_addr[16]));
 sky130_fd_sc_hd__clkbuf_2 output142 (.A(net142),
    .X(mem_addr[17]));
 sky130_fd_sc_hd__clkbuf_2 output143 (.A(net143),
    .X(mem_addr[18]));
 sky130_fd_sc_hd__clkbuf_2 output144 (.A(net144),
    .X(mem_addr[19]));
 sky130_fd_sc_hd__clkbuf_2 output145 (.A(net145),
    .X(mem_addr[1]));
 sky130_fd_sc_hd__clkbuf_2 output146 (.A(net146),
    .X(mem_addr[20]));
 sky130_fd_sc_hd__clkbuf_2 output147 (.A(net147),
    .X(mem_addr[21]));
 sky130_fd_sc_hd__clkbuf_2 output148 (.A(net148),
    .X(mem_addr[22]));
 sky130_fd_sc_hd__clkbuf_2 output149 (.A(net149),
    .X(mem_addr[23]));
 sky130_fd_sc_hd__clkbuf_2 output150 (.A(net150),
    .X(mem_addr[24]));
 sky130_fd_sc_hd__clkbuf_2 output151 (.A(net151),
    .X(mem_addr[25]));
 sky130_fd_sc_hd__clkbuf_2 output152 (.A(net152),
    .X(mem_addr[26]));
 sky130_fd_sc_hd__clkbuf_2 output153 (.A(net153),
    .X(mem_addr[27]));
 sky130_fd_sc_hd__clkbuf_2 output154 (.A(net154),
    .X(mem_addr[28]));
 sky130_fd_sc_hd__clkbuf_2 output155 (.A(net155),
    .X(mem_addr[29]));
 sky130_fd_sc_hd__clkbuf_2 output156 (.A(net156),
    .X(mem_addr[2]));
 sky130_fd_sc_hd__clkbuf_2 output157 (.A(net157),
    .X(mem_addr[30]));
 sky130_fd_sc_hd__clkbuf_2 output158 (.A(net158),
    .X(mem_addr[31]));
 sky130_fd_sc_hd__clkbuf_2 output159 (.A(net159),
    .X(mem_addr[3]));
 sky130_fd_sc_hd__clkbuf_2 output160 (.A(net160),
    .X(mem_addr[4]));
 sky130_fd_sc_hd__clkbuf_2 output161 (.A(net161),
    .X(mem_addr[5]));
 sky130_fd_sc_hd__clkbuf_2 output162 (.A(net162),
    .X(mem_addr[6]));
 sky130_fd_sc_hd__clkbuf_2 output163 (.A(net163),
    .X(mem_addr[7]));
 sky130_fd_sc_hd__clkbuf_2 output164 (.A(net164),
    .X(mem_addr[8]));
 sky130_fd_sc_hd__clkbuf_2 output165 (.A(net165),
    .X(mem_addr[9]));
 sky130_fd_sc_hd__clkbuf_2 output166 (.A(net166),
    .X(mem_instr));
 sky130_fd_sc_hd__clkbuf_2 output167 (.A(net167),
    .X(mem_la_addr[0]));
 sky130_fd_sc_hd__clkbuf_2 output168 (.A(net168),
    .X(mem_la_addr[10]));
 sky130_fd_sc_hd__clkbuf_2 output169 (.A(net169),
    .X(mem_la_addr[11]));
 sky130_fd_sc_hd__clkbuf_2 output170 (.A(net170),
    .X(mem_la_addr[12]));
 sky130_fd_sc_hd__clkbuf_2 output171 (.A(net171),
    .X(mem_la_addr[13]));
 sky130_fd_sc_hd__clkbuf_2 output172 (.A(net172),
    .X(mem_la_addr[14]));
 sky130_fd_sc_hd__clkbuf_2 output173 (.A(net173),
    .X(mem_la_addr[15]));
 sky130_fd_sc_hd__clkbuf_2 output174 (.A(net174),
    .X(mem_la_addr[16]));
 sky130_fd_sc_hd__clkbuf_2 output175 (.A(net175),
    .X(mem_la_addr[17]));
 sky130_fd_sc_hd__clkbuf_2 output176 (.A(net176),
    .X(mem_la_addr[18]));
 sky130_fd_sc_hd__clkbuf_2 output177 (.A(net177),
    .X(mem_la_addr[19]));
 sky130_fd_sc_hd__clkbuf_2 output178 (.A(net178),
    .X(mem_la_addr[1]));
 sky130_fd_sc_hd__clkbuf_2 output179 (.A(net179),
    .X(mem_la_addr[20]));
 sky130_fd_sc_hd__clkbuf_2 output180 (.A(net180),
    .X(mem_la_addr[21]));
 sky130_fd_sc_hd__clkbuf_2 output181 (.A(net181),
    .X(mem_la_addr[22]));
 sky130_fd_sc_hd__clkbuf_2 output182 (.A(net182),
    .X(mem_la_addr[23]));
 sky130_fd_sc_hd__clkbuf_2 output183 (.A(net183),
    .X(mem_la_addr[24]));
 sky130_fd_sc_hd__clkbuf_2 output184 (.A(net184),
    .X(mem_la_addr[25]));
 sky130_fd_sc_hd__clkbuf_2 output185 (.A(net185),
    .X(mem_la_addr[26]));
 sky130_fd_sc_hd__clkbuf_2 output186 (.A(net186),
    .X(mem_la_addr[27]));
 sky130_fd_sc_hd__clkbuf_2 output187 (.A(net187),
    .X(mem_la_addr[28]));
 sky130_fd_sc_hd__clkbuf_2 output188 (.A(net188),
    .X(mem_la_addr[29]));
 sky130_fd_sc_hd__clkbuf_2 output189 (.A(net189),
    .X(mem_la_addr[2]));
 sky130_fd_sc_hd__clkbuf_2 output190 (.A(net190),
    .X(mem_la_addr[30]));
 sky130_fd_sc_hd__clkbuf_2 output191 (.A(net191),
    .X(mem_la_addr[31]));
 sky130_fd_sc_hd__clkbuf_2 output192 (.A(net192),
    .X(mem_la_addr[3]));
 sky130_fd_sc_hd__clkbuf_2 output193 (.A(net193),
    .X(mem_la_addr[4]));
 sky130_fd_sc_hd__clkbuf_2 output194 (.A(net194),
    .X(mem_la_addr[5]));
 sky130_fd_sc_hd__clkbuf_2 output195 (.A(net195),
    .X(mem_la_addr[6]));
 sky130_fd_sc_hd__clkbuf_2 output196 (.A(net196),
    .X(mem_la_addr[7]));
 sky130_fd_sc_hd__clkbuf_2 output197 (.A(net197),
    .X(mem_la_addr[8]));
 sky130_fd_sc_hd__clkbuf_2 output198 (.A(net198),
    .X(mem_la_addr[9]));
 sky130_fd_sc_hd__clkbuf_2 output199 (.A(net199),
    .X(mem_la_read));
 sky130_fd_sc_hd__clkbuf_2 output200 (.A(net506),
    .X(mem_la_wdata[0]));
 sky130_fd_sc_hd__clkbuf_2 output201 (.A(net201),
    .X(mem_la_wdata[10]));
 sky130_fd_sc_hd__clkbuf_2 output202 (.A(net202),
    .X(mem_la_wdata[11]));
 sky130_fd_sc_hd__clkbuf_2 output203 (.A(net203),
    .X(mem_la_wdata[12]));
 sky130_fd_sc_hd__clkbuf_2 output204 (.A(net204),
    .X(mem_la_wdata[13]));
 sky130_fd_sc_hd__clkbuf_2 output205 (.A(net205),
    .X(mem_la_wdata[14]));
 sky130_fd_sc_hd__clkbuf_2 output206 (.A(net206),
    .X(mem_la_wdata[15]));
 sky130_fd_sc_hd__clkbuf_2 output207 (.A(net207),
    .X(mem_la_wdata[16]));
 sky130_fd_sc_hd__clkbuf_2 output208 (.A(net208),
    .X(mem_la_wdata[17]));
 sky130_fd_sc_hd__clkbuf_2 output209 (.A(net209),
    .X(mem_la_wdata[18]));
 sky130_fd_sc_hd__clkbuf_2 output210 (.A(net210),
    .X(mem_la_wdata[19]));
 sky130_fd_sc_hd__clkbuf_2 output211 (.A(net211),
    .X(mem_la_wdata[1]));
 sky130_fd_sc_hd__clkbuf_2 output212 (.A(net212),
    .X(mem_la_wdata[20]));
 sky130_fd_sc_hd__clkbuf_2 output213 (.A(net213),
    .X(mem_la_wdata[21]));
 sky130_fd_sc_hd__clkbuf_2 output214 (.A(net214),
    .X(mem_la_wdata[22]));
 sky130_fd_sc_hd__clkbuf_2 output215 (.A(net215),
    .X(mem_la_wdata[23]));
 sky130_fd_sc_hd__clkbuf_2 output216 (.A(net216),
    .X(mem_la_wdata[24]));
 sky130_fd_sc_hd__clkbuf_2 output217 (.A(net217),
    .X(mem_la_wdata[25]));
 sky130_fd_sc_hd__clkbuf_2 output218 (.A(net218),
    .X(mem_la_wdata[26]));
 sky130_fd_sc_hd__clkbuf_2 output219 (.A(net219),
    .X(mem_la_wdata[27]));
 sky130_fd_sc_hd__clkbuf_2 output220 (.A(net220),
    .X(mem_la_wdata[28]));
 sky130_fd_sc_hd__clkbuf_2 output221 (.A(net221),
    .X(mem_la_wdata[29]));
 sky130_fd_sc_hd__clkbuf_2 output222 (.A(net504),
    .X(mem_la_wdata[2]));
 sky130_fd_sc_hd__clkbuf_2 output223 (.A(net223),
    .X(mem_la_wdata[30]));
 sky130_fd_sc_hd__clkbuf_2 output224 (.A(net224),
    .X(mem_la_wdata[31]));
 sky130_fd_sc_hd__clkbuf_2 output225 (.A(net225),
    .X(mem_la_wdata[3]));
 sky130_fd_sc_hd__clkbuf_2 output226 (.A(net226),
    .X(mem_la_wdata[4]));
 sky130_fd_sc_hd__clkbuf_2 output227 (.A(net227),
    .X(mem_la_wdata[5]));
 sky130_fd_sc_hd__clkbuf_2 output228 (.A(net228),
    .X(mem_la_wdata[6]));
 sky130_fd_sc_hd__clkbuf_2 output229 (.A(net229),
    .X(mem_la_wdata[7]));
 sky130_fd_sc_hd__clkbuf_2 output230 (.A(net230),
    .X(mem_la_wdata[8]));
 sky130_fd_sc_hd__clkbuf_2 output231 (.A(net231),
    .X(mem_la_wdata[9]));
 sky130_fd_sc_hd__clkbuf_2 output232 (.A(net232),
    .X(mem_la_write));
 sky130_fd_sc_hd__clkbuf_2 output233 (.A(net233),
    .X(mem_la_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_2 output234 (.A(net234),
    .X(mem_la_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_2 output235 (.A(net235),
    .X(mem_la_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_2 output236 (.A(net236),
    .X(mem_la_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_2 output237 (.A(net237),
    .X(mem_valid));
 sky130_fd_sc_hd__clkbuf_2 output238 (.A(net238),
    .X(mem_wdata[0]));
 sky130_fd_sc_hd__clkbuf_2 output239 (.A(net239),
    .X(mem_wdata[10]));
 sky130_fd_sc_hd__clkbuf_2 output240 (.A(net240),
    .X(mem_wdata[11]));
 sky130_fd_sc_hd__clkbuf_2 output241 (.A(net241),
    .X(mem_wdata[12]));
 sky130_fd_sc_hd__clkbuf_2 output242 (.A(net242),
    .X(mem_wdata[13]));
 sky130_fd_sc_hd__clkbuf_2 output243 (.A(net243),
    .X(mem_wdata[14]));
 sky130_fd_sc_hd__clkbuf_2 output244 (.A(net244),
    .X(mem_wdata[15]));
 sky130_fd_sc_hd__clkbuf_2 output245 (.A(net245),
    .X(mem_wdata[16]));
 sky130_fd_sc_hd__clkbuf_2 output246 (.A(net246),
    .X(mem_wdata[17]));
 sky130_fd_sc_hd__clkbuf_2 output247 (.A(net247),
    .X(mem_wdata[18]));
 sky130_fd_sc_hd__clkbuf_2 output248 (.A(net248),
    .X(mem_wdata[19]));
 sky130_fd_sc_hd__clkbuf_2 output249 (.A(net249),
    .X(mem_wdata[1]));
 sky130_fd_sc_hd__clkbuf_2 output250 (.A(net250),
    .X(mem_wdata[20]));
 sky130_fd_sc_hd__clkbuf_2 output251 (.A(net251),
    .X(mem_wdata[21]));
 sky130_fd_sc_hd__clkbuf_2 output252 (.A(net252),
    .X(mem_wdata[22]));
 sky130_fd_sc_hd__clkbuf_2 output253 (.A(net253),
    .X(mem_wdata[23]));
 sky130_fd_sc_hd__clkbuf_2 output254 (.A(net254),
    .X(mem_wdata[24]));
 sky130_fd_sc_hd__clkbuf_2 output255 (.A(net255),
    .X(mem_wdata[25]));
 sky130_fd_sc_hd__clkbuf_2 output256 (.A(net256),
    .X(mem_wdata[26]));
 sky130_fd_sc_hd__clkbuf_2 output257 (.A(net257),
    .X(mem_wdata[27]));
 sky130_fd_sc_hd__clkbuf_2 output258 (.A(net258),
    .X(mem_wdata[28]));
 sky130_fd_sc_hd__clkbuf_2 output259 (.A(net259),
    .X(mem_wdata[29]));
 sky130_fd_sc_hd__clkbuf_2 output260 (.A(net260),
    .X(mem_wdata[2]));
 sky130_fd_sc_hd__clkbuf_2 output261 (.A(net261),
    .X(mem_wdata[30]));
 sky130_fd_sc_hd__clkbuf_2 output262 (.A(net262),
    .X(mem_wdata[31]));
 sky130_fd_sc_hd__clkbuf_2 output263 (.A(net263),
    .X(mem_wdata[3]));
 sky130_fd_sc_hd__clkbuf_2 output264 (.A(net264),
    .X(mem_wdata[4]));
 sky130_fd_sc_hd__clkbuf_2 output265 (.A(net265),
    .X(mem_wdata[5]));
 sky130_fd_sc_hd__clkbuf_2 output266 (.A(net266),
    .X(mem_wdata[6]));
 sky130_fd_sc_hd__clkbuf_2 output267 (.A(net267),
    .X(mem_wdata[7]));
 sky130_fd_sc_hd__clkbuf_2 output268 (.A(net268),
    .X(mem_wdata[8]));
 sky130_fd_sc_hd__clkbuf_2 output269 (.A(net269),
    .X(mem_wdata[9]));
 sky130_fd_sc_hd__clkbuf_2 output270 (.A(net270),
    .X(mem_wstrb[0]));
 sky130_fd_sc_hd__clkbuf_2 output271 (.A(net271),
    .X(mem_wstrb[1]));
 sky130_fd_sc_hd__clkbuf_2 output272 (.A(net272),
    .X(mem_wstrb[2]));
 sky130_fd_sc_hd__clkbuf_2 output273 (.A(net273),
    .X(mem_wstrb[3]));
 sky130_fd_sc_hd__clkbuf_2 output274 (.A(net274),
    .X(pcpi_insn[0]));
 sky130_fd_sc_hd__clkbuf_2 output275 (.A(net275),
    .X(pcpi_insn[10]));
 sky130_fd_sc_hd__clkbuf_2 output276 (.A(net276),
    .X(pcpi_insn[11]));
 sky130_fd_sc_hd__clkbuf_2 output277 (.A(net277),
    .X(pcpi_insn[12]));
 sky130_fd_sc_hd__clkbuf_2 output278 (.A(net278),
    .X(pcpi_insn[13]));
 sky130_fd_sc_hd__clkbuf_2 output279 (.A(net279),
    .X(pcpi_insn[14]));
 sky130_fd_sc_hd__clkbuf_2 output280 (.A(net280),
    .X(pcpi_insn[15]));
 sky130_fd_sc_hd__clkbuf_2 output281 (.A(net281),
    .X(pcpi_insn[16]));
 sky130_fd_sc_hd__clkbuf_2 output282 (.A(net282),
    .X(pcpi_insn[17]));
 sky130_fd_sc_hd__clkbuf_2 output283 (.A(net283),
    .X(pcpi_insn[18]));
 sky130_fd_sc_hd__clkbuf_2 output284 (.A(net284),
    .X(pcpi_insn[19]));
 sky130_fd_sc_hd__clkbuf_2 output285 (.A(net285),
    .X(pcpi_insn[1]));
 sky130_fd_sc_hd__clkbuf_2 output286 (.A(net286),
    .X(pcpi_insn[20]));
 sky130_fd_sc_hd__clkbuf_2 output287 (.A(net287),
    .X(pcpi_insn[21]));
 sky130_fd_sc_hd__clkbuf_2 output288 (.A(net288),
    .X(pcpi_insn[22]));
 sky130_fd_sc_hd__clkbuf_2 output289 (.A(net289),
    .X(pcpi_insn[23]));
 sky130_fd_sc_hd__clkbuf_2 output290 (.A(net290),
    .X(pcpi_insn[24]));
 sky130_fd_sc_hd__clkbuf_2 output291 (.A(net291),
    .X(pcpi_insn[25]));
 sky130_fd_sc_hd__clkbuf_2 output292 (.A(net292),
    .X(pcpi_insn[26]));
 sky130_fd_sc_hd__clkbuf_2 output293 (.A(net293),
    .X(pcpi_insn[27]));
 sky130_fd_sc_hd__clkbuf_2 output294 (.A(net294),
    .X(pcpi_insn[28]));
 sky130_fd_sc_hd__clkbuf_2 output295 (.A(net295),
    .X(pcpi_insn[29]));
 sky130_fd_sc_hd__clkbuf_2 output296 (.A(net296),
    .X(pcpi_insn[2]));
 sky130_fd_sc_hd__clkbuf_2 output297 (.A(net297),
    .X(pcpi_insn[30]));
 sky130_fd_sc_hd__clkbuf_2 output298 (.A(net298),
    .X(pcpi_insn[31]));
 sky130_fd_sc_hd__clkbuf_2 output299 (.A(net299),
    .X(pcpi_insn[3]));
 sky130_fd_sc_hd__clkbuf_2 output300 (.A(net300),
    .X(pcpi_insn[4]));
 sky130_fd_sc_hd__clkbuf_2 output301 (.A(net301),
    .X(pcpi_insn[5]));
 sky130_fd_sc_hd__clkbuf_2 output302 (.A(net302),
    .X(pcpi_insn[6]));
 sky130_fd_sc_hd__clkbuf_2 output303 (.A(net303),
    .X(pcpi_insn[7]));
 sky130_fd_sc_hd__clkbuf_2 output304 (.A(net304),
    .X(pcpi_insn[8]));
 sky130_fd_sc_hd__clkbuf_2 output305 (.A(net305),
    .X(pcpi_insn[9]));
 sky130_fd_sc_hd__clkbuf_2 output306 (.A(net306),
    .X(pcpi_rs1[0]));
 sky130_fd_sc_hd__clkbuf_2 output307 (.A(net307),
    .X(pcpi_rs1[10]));
 sky130_fd_sc_hd__clkbuf_2 output308 (.A(net308),
    .X(pcpi_rs1[11]));
 sky130_fd_sc_hd__clkbuf_2 output309 (.A(net309),
    .X(pcpi_rs1[12]));
 sky130_fd_sc_hd__clkbuf_2 output310 (.A(net310),
    .X(pcpi_rs1[13]));
 sky130_fd_sc_hd__clkbuf_2 output311 (.A(net311),
    .X(pcpi_rs1[14]));
 sky130_fd_sc_hd__clkbuf_2 output312 (.A(net312),
    .X(pcpi_rs1[15]));
 sky130_fd_sc_hd__clkbuf_2 output313 (.A(net313),
    .X(pcpi_rs1[16]));
 sky130_fd_sc_hd__clkbuf_2 output314 (.A(net314),
    .X(pcpi_rs1[17]));
 sky130_fd_sc_hd__clkbuf_2 output315 (.A(net315),
    .X(pcpi_rs1[18]));
 sky130_fd_sc_hd__clkbuf_2 output316 (.A(net316),
    .X(pcpi_rs1[19]));
 sky130_fd_sc_hd__clkbuf_2 output317 (.A(net317),
    .X(pcpi_rs1[1]));
 sky130_fd_sc_hd__clkbuf_2 output318 (.A(net318),
    .X(pcpi_rs1[20]));
 sky130_fd_sc_hd__clkbuf_2 output319 (.A(net319),
    .X(pcpi_rs1[21]));
 sky130_fd_sc_hd__clkbuf_2 output320 (.A(net320),
    .X(pcpi_rs1[22]));
 sky130_fd_sc_hd__clkbuf_2 output321 (.A(net321),
    .X(pcpi_rs1[23]));
 sky130_fd_sc_hd__clkbuf_2 output322 (.A(net322),
    .X(pcpi_rs1[24]));
 sky130_fd_sc_hd__clkbuf_2 output323 (.A(net323),
    .X(pcpi_rs1[25]));
 sky130_fd_sc_hd__clkbuf_2 output324 (.A(net324),
    .X(pcpi_rs1[26]));
 sky130_fd_sc_hd__clkbuf_2 output325 (.A(net325),
    .X(pcpi_rs1[27]));
 sky130_fd_sc_hd__clkbuf_2 output326 (.A(net326),
    .X(pcpi_rs1[28]));
 sky130_fd_sc_hd__clkbuf_2 output327 (.A(net327),
    .X(pcpi_rs1[29]));
 sky130_fd_sc_hd__clkbuf_2 output328 (.A(net328),
    .X(pcpi_rs1[2]));
 sky130_fd_sc_hd__clkbuf_2 output329 (.A(net329),
    .X(pcpi_rs1[30]));
 sky130_fd_sc_hd__clkbuf_2 output330 (.A(net330),
    .X(pcpi_rs1[31]));
 sky130_fd_sc_hd__clkbuf_2 output331 (.A(net331),
    .X(pcpi_rs1[3]));
 sky130_fd_sc_hd__clkbuf_2 output332 (.A(net332),
    .X(pcpi_rs1[4]));
 sky130_fd_sc_hd__clkbuf_2 output333 (.A(net333),
    .X(pcpi_rs1[5]));
 sky130_fd_sc_hd__clkbuf_2 output334 (.A(net334),
    .X(pcpi_rs1[6]));
 sky130_fd_sc_hd__clkbuf_2 output335 (.A(net335),
    .X(pcpi_rs1[7]));
 sky130_fd_sc_hd__clkbuf_2 output336 (.A(net336),
    .X(pcpi_rs1[8]));
 sky130_fd_sc_hd__clkbuf_2 output337 (.A(net337),
    .X(pcpi_rs1[9]));
 sky130_fd_sc_hd__clkbuf_2 output338 (.A(net338),
    .X(pcpi_rs2[0]));
 sky130_fd_sc_hd__clkbuf_2 output339 (.A(net339),
    .X(pcpi_rs2[10]));
 sky130_fd_sc_hd__clkbuf_2 output340 (.A(net340),
    .X(pcpi_rs2[11]));
 sky130_fd_sc_hd__clkbuf_2 output341 (.A(net341),
    .X(pcpi_rs2[12]));
 sky130_fd_sc_hd__clkbuf_2 output342 (.A(net342),
    .X(pcpi_rs2[13]));
 sky130_fd_sc_hd__clkbuf_2 output343 (.A(net343),
    .X(pcpi_rs2[14]));
 sky130_fd_sc_hd__clkbuf_2 output344 (.A(net344),
    .X(pcpi_rs2[15]));
 sky130_fd_sc_hd__clkbuf_2 output345 (.A(net345),
    .X(pcpi_rs2[16]));
 sky130_fd_sc_hd__clkbuf_2 output346 (.A(net346),
    .X(pcpi_rs2[17]));
 sky130_fd_sc_hd__clkbuf_2 output347 (.A(net347),
    .X(pcpi_rs2[18]));
 sky130_fd_sc_hd__clkbuf_2 output348 (.A(net348),
    .X(pcpi_rs2[19]));
 sky130_fd_sc_hd__clkbuf_2 output349 (.A(net349),
    .X(pcpi_rs2[1]));
 sky130_fd_sc_hd__clkbuf_2 output350 (.A(net350),
    .X(pcpi_rs2[20]));
 sky130_fd_sc_hd__clkbuf_2 output351 (.A(net351),
    .X(pcpi_rs2[21]));
 sky130_fd_sc_hd__clkbuf_2 output352 (.A(net352),
    .X(pcpi_rs2[22]));
 sky130_fd_sc_hd__clkbuf_2 output353 (.A(net353),
    .X(pcpi_rs2[23]));
 sky130_fd_sc_hd__clkbuf_2 output354 (.A(net354),
    .X(pcpi_rs2[24]));
 sky130_fd_sc_hd__clkbuf_2 output355 (.A(net355),
    .X(pcpi_rs2[25]));
 sky130_fd_sc_hd__clkbuf_2 output356 (.A(net356),
    .X(pcpi_rs2[26]));
 sky130_fd_sc_hd__clkbuf_2 output357 (.A(net357),
    .X(pcpi_rs2[27]));
 sky130_fd_sc_hd__clkbuf_2 output358 (.A(net358),
    .X(pcpi_rs2[28]));
 sky130_fd_sc_hd__clkbuf_2 output359 (.A(net359),
    .X(pcpi_rs2[29]));
 sky130_fd_sc_hd__clkbuf_2 output360 (.A(net360),
    .X(pcpi_rs2[2]));
 sky130_fd_sc_hd__clkbuf_2 output361 (.A(net361),
    .X(pcpi_rs2[30]));
 sky130_fd_sc_hd__clkbuf_2 output362 (.A(net362),
    .X(pcpi_rs2[31]));
 sky130_fd_sc_hd__clkbuf_2 output363 (.A(net363),
    .X(pcpi_rs2[3]));
 sky130_fd_sc_hd__clkbuf_2 output364 (.A(net364),
    .X(pcpi_rs2[4]));
 sky130_fd_sc_hd__clkbuf_2 output365 (.A(net365),
    .X(pcpi_rs2[5]));
 sky130_fd_sc_hd__clkbuf_2 output366 (.A(net366),
    .X(pcpi_rs2[6]));
 sky130_fd_sc_hd__clkbuf_2 output367 (.A(net367),
    .X(pcpi_rs2[7]));
 sky130_fd_sc_hd__clkbuf_2 output368 (.A(net368),
    .X(pcpi_rs2[8]));
 sky130_fd_sc_hd__clkbuf_2 output369 (.A(net369),
    .X(pcpi_rs2[9]));
 sky130_fd_sc_hd__clkbuf_2 output370 (.A(net370),
    .X(pcpi_valid));
 sky130_fd_sc_hd__clkbuf_2 output371 (.A(net371),
    .X(trace_data[0]));
 sky130_fd_sc_hd__clkbuf_2 output372 (.A(net372),
    .X(trace_data[10]));
 sky130_fd_sc_hd__clkbuf_2 output373 (.A(net373),
    .X(trace_data[11]));
 sky130_fd_sc_hd__clkbuf_2 output374 (.A(net374),
    .X(trace_data[12]));
 sky130_fd_sc_hd__clkbuf_2 output375 (.A(net375),
    .X(trace_data[13]));
 sky130_fd_sc_hd__clkbuf_2 output376 (.A(net376),
    .X(trace_data[14]));
 sky130_fd_sc_hd__clkbuf_2 output377 (.A(net377),
    .X(trace_data[15]));
 sky130_fd_sc_hd__clkbuf_2 output378 (.A(net378),
    .X(trace_data[16]));
 sky130_fd_sc_hd__clkbuf_2 output379 (.A(net379),
    .X(trace_data[17]));
 sky130_fd_sc_hd__clkbuf_2 output380 (.A(net380),
    .X(trace_data[18]));
 sky130_fd_sc_hd__clkbuf_2 output381 (.A(net381),
    .X(trace_data[19]));
 sky130_fd_sc_hd__clkbuf_2 output382 (.A(net382),
    .X(trace_data[1]));
 sky130_fd_sc_hd__clkbuf_2 output383 (.A(net383),
    .X(trace_data[20]));
 sky130_fd_sc_hd__clkbuf_2 output384 (.A(net384),
    .X(trace_data[21]));
 sky130_fd_sc_hd__clkbuf_2 output385 (.A(net385),
    .X(trace_data[22]));
 sky130_fd_sc_hd__clkbuf_2 output386 (.A(net386),
    .X(trace_data[23]));
 sky130_fd_sc_hd__clkbuf_2 output387 (.A(net387),
    .X(trace_data[24]));
 sky130_fd_sc_hd__clkbuf_2 output388 (.A(net388),
    .X(trace_data[25]));
 sky130_fd_sc_hd__clkbuf_2 output389 (.A(net389),
    .X(trace_data[26]));
 sky130_fd_sc_hd__clkbuf_2 output390 (.A(net390),
    .X(trace_data[27]));
 sky130_fd_sc_hd__clkbuf_2 output391 (.A(net391),
    .X(trace_data[28]));
 sky130_fd_sc_hd__clkbuf_2 output392 (.A(net392),
    .X(trace_data[29]));
 sky130_fd_sc_hd__clkbuf_2 output393 (.A(net393),
    .X(trace_data[2]));
 sky130_fd_sc_hd__clkbuf_2 output394 (.A(net394),
    .X(trace_data[30]));
 sky130_fd_sc_hd__clkbuf_2 output395 (.A(net395),
    .X(trace_data[31]));
 sky130_fd_sc_hd__clkbuf_2 output396 (.A(net396),
    .X(trace_data[32]));
 sky130_fd_sc_hd__clkbuf_2 output397 (.A(net397),
    .X(trace_data[33]));
 sky130_fd_sc_hd__clkbuf_2 output398 (.A(net398),
    .X(trace_data[34]));
 sky130_fd_sc_hd__clkbuf_2 output399 (.A(net399),
    .X(trace_data[35]));
 sky130_fd_sc_hd__clkbuf_2 output400 (.A(net400),
    .X(trace_data[3]));
 sky130_fd_sc_hd__clkbuf_2 output401 (.A(net401),
    .X(trace_data[4]));
 sky130_fd_sc_hd__clkbuf_2 output402 (.A(net402),
    .X(trace_data[5]));
 sky130_fd_sc_hd__clkbuf_2 output403 (.A(net403),
    .X(trace_data[6]));
 sky130_fd_sc_hd__clkbuf_2 output404 (.A(net404),
    .X(trace_data[7]));
 sky130_fd_sc_hd__clkbuf_2 output405 (.A(net405),
    .X(trace_data[8]));
 sky130_fd_sc_hd__clkbuf_2 output406 (.A(net406),
    .X(trace_data[9]));
 sky130_fd_sc_hd__clkbuf_2 output407 (.A(net407),
    .X(trace_valid));
 sky130_fd_sc_hd__clkbuf_2 output408 (.A(net408),
    .X(trap));
 sky130_fd_sc_hd__buf_12 repeater409 (.A(_11327_),
    .X(net409));
 sky130_fd_sc_hd__buf_6 repeater410 (.A(_14332_),
    .X(net410));
 sky130_fd_sc_hd__buf_6 repeater411 (.A(_13720_),
    .X(net411));
 sky130_fd_sc_hd__buf_8 repeater412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__buf_8 repeater413 (.A(_00308_),
    .X(net413));
 sky130_fd_sc_hd__buf_8 repeater414 (.A(_19824_),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_8 repeater415 (.A(_19823_),
    .X(net415));
 sky130_fd_sc_hd__buf_8 repeater416 (.A(_19822_),
    .X(net416));
 sky130_fd_sc_hd__buf_8 repeater417 (.A(_19821_),
    .X(net417));
 sky130_fd_sc_hd__buf_6 repeater418 (.A(_19479_),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_8 repeater419 (.A(_19478_),
    .X(net419));
 sky130_fd_sc_hd__buf_8 repeater420 (.A(_19477_),
    .X(net420));
 sky130_fd_sc_hd__buf_4 repeater421 (.A(_19476_),
    .X(net421));
 sky130_fd_sc_hd__buf_8 repeater422 (.A(_18635_),
    .X(net422));
 sky130_fd_sc_hd__buf_8 repeater423 (.A(_19480_),
    .X(net423));
 sky130_fd_sc_hd__buf_12 repeater424 (.A(_02217_),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_8 repeater425 (.A(_18600_),
    .X(net425));
 sky130_fd_sc_hd__buf_8 repeater426 (.A(_18581_),
    .X(net426));
 sky130_fd_sc_hd__buf_6 repeater427 (.A(_18580_),
    .X(net427));
 sky130_fd_sc_hd__buf_12 repeater428 (.A(_20894_),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_8 repeater429 (.A(_02069_),
    .X(net429));
 sky130_fd_sc_hd__buf_4 repeater430 (.A(_02069_),
    .X(net430));
 sky130_fd_sc_hd__buf_8 repeater431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_8 repeater432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_8 repeater433 (.A(_01683_),
    .X(net433));
 sky130_fd_sc_hd__buf_4 repeater434 (.A(_01683_),
    .X(net434));
 sky130_fd_sc_hd__buf_8 repeater435 (.A(_19889_),
    .X(net435));
 sky130_fd_sc_hd__buf_8 repeater436 (.A(_18606_),
    .X(net436));
 sky130_fd_sc_hd__buf_8 repeater437 (.A(_18565_),
    .X(net437));
 sky130_fd_sc_hd__buf_8 repeater438 (.A(_08745_),
    .X(net438));
 sky130_fd_sc_hd__buf_6 repeater439 (.A(_08044_),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_8 repeater440 (.A(_07289_),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_8 repeater441 (.A(_06929_),
    .X(net441));
 sky130_fd_sc_hd__buf_8 repeater442 (.A(_06829_),
    .X(net442));
 sky130_fd_sc_hd__buf_6 repeater443 (.A(_06460_),
    .X(net443));
 sky130_fd_sc_hd__buf_8 repeater444 (.A(_06434_),
    .X(net444));
 sky130_fd_sc_hd__buf_6 repeater445 (.A(_06352_),
    .X(net445));
 sky130_fd_sc_hd__buf_6 repeater446 (.A(_06263_),
    .X(net446));
 sky130_fd_sc_hd__buf_8 repeater447 (.A(_05803_),
    .X(net447));
 sky130_fd_sc_hd__buf_4 repeater448 (.A(_05737_),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_8 repeater449 (.A(_05669_),
    .X(net449));
 sky130_fd_sc_hd__buf_8 repeater450 (.A(_05616_),
    .X(net450));
 sky130_fd_sc_hd__buf_4 repeater451 (.A(_05551_),
    .X(net451));
 sky130_fd_sc_hd__buf_6 repeater452 (.A(_05279_),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_8 repeater453 (.A(_04841_),
    .X(net453));
 sky130_fd_sc_hd__buf_6 repeater454 (.A(_19882_),
    .X(net454));
 sky130_fd_sc_hd__buf_6 repeater455 (.A(_19671_),
    .X(net455));
 sky130_fd_sc_hd__buf_8 repeater456 (.A(_19660_),
    .X(net456));
 sky130_fd_sc_hd__buf_4 repeater457 (.A(_19656_),
    .X(net457));
 sky130_fd_sc_hd__buf_6 repeater458 (.A(_19642_),
    .X(net458));
 sky130_fd_sc_hd__buf_8 repeater459 (.A(net462),
    .X(net459));
 sky130_fd_sc_hd__buf_8 repeater460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_8 repeater461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_8 repeater462 (.A(_00301_),
    .X(net462));
 sky130_fd_sc_hd__buf_4 repeater463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_8 repeater464 (.A(_01706_),
    .X(net464));
 sky130_fd_sc_hd__buf_6 repeater465 (.A(_18469_),
    .X(net465));
 sky130_fd_sc_hd__buf_12 repeater466 (.A(_00368_),
    .X(net466));
 sky130_fd_sc_hd__buf_12 repeater467 (.A(_00368_),
    .X(net467));
 sky130_fd_sc_hd__buf_8 repeater468 (.A(_13118_),
    .X(net468));
 sky130_fd_sc_hd__buf_6 repeater469 (.A(_10836_),
    .X(net469));
 sky130_fd_sc_hd__buf_6 repeater470 (.A(_07561_),
    .X(net470));
 sky130_fd_sc_hd__buf_6 repeater471 (.A(_07042_),
    .X(net471));
 sky130_fd_sc_hd__buf_4 repeater472 (.A(_06215_),
    .X(net472));
 sky130_fd_sc_hd__buf_6 repeater473 (.A(_06031_),
    .X(net473));
 sky130_fd_sc_hd__buf_8 repeater474 (.A(_04839_),
    .X(net474));
 sky130_fd_sc_hd__buf_8 repeater475 (.A(_01304_),
    .X(net475));
 sky130_fd_sc_hd__buf_8 repeater476 (.A(_19686_),
    .X(net476));
 sky130_fd_sc_hd__buf_8 repeater477 (.A(_19652_),
    .X(net477));
 sky130_fd_sc_hd__buf_6 repeater478 (.A(_19650_),
    .X(net478));
 sky130_fd_sc_hd__buf_12 repeater479 (.A(mem_xfer),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_16 repeater480 (.A(_00357_),
    .X(net480));
 sky130_fd_sc_hd__buf_12 repeater481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_12 repeater482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_12 repeater483 (.A(net488),
    .X(net483));
 sky130_fd_sc_hd__buf_12 repeater484 (.A(net485),
    .X(net484));
 sky130_fd_sc_hd__buf_12 repeater485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__buf_12 repeater486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__buf_8 repeater487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_12 repeater488 (.A(_00358_),
    .X(net488));
 sky130_fd_sc_hd__buf_12 repeater489 (.A(net491),
    .X(net489));
 sky130_fd_sc_hd__buf_12 repeater490 (.A(net491),
    .X(net490));
 sky130_fd_sc_hd__buf_12 repeater491 (.A(_00360_),
    .X(net491));
 sky130_fd_sc_hd__buf_12 repeater492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_12 repeater493 (.A(_00362_),
    .X(net493));
 sky130_fd_sc_hd__buf_6 repeater494 (.A(_11094_),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_8 repeater495 (.A(_05207_),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_8 repeater496 (.A(_01816_),
    .X(net496));
 sky130_fd_sc_hd__buf_4 repeater497 (.A(_19880_),
    .X(net497));
 sky130_fd_sc_hd__buf_8 repeater498 (.A(_19579_),
    .X(net498));
 sky130_fd_sc_hd__buf_8 repeater499 (.A(_19447_),
    .X(net499));
 sky130_fd_sc_hd__buf_8 repeater500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__buf_8 repeater501 (.A(_00297_),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_16 repeater502 (.A(net226),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_16 repeater503 (.A(net225),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_16 repeater504 (.A(net222),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_16 repeater505 (.A(net211),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_16 repeater506 (.A(net200),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_16 repeater507 (.A(\cpu_state[3] ),
    .X(net507));
 sky130_fd_sc_hd__buf_12 repeater508 (.A(\cpu_state[2] ),
    .X(net508));
 sky130_fd_sc_hd__clkbuf_16 repeater509 (.A(\pcpi_mul.shift_out ),
    .X(net509));
 sky130_fd_sc_hd__buf_8 repeater510 (.A(net7),
    .X(net510));
 sky130_fd_sc_hd__buf_8 repeater511 (.A(net65),
    .X(net511));
 sky130_fd_sc_hd__buf_8 repeater512 (.A(net60),
    .X(net512));
 sky130_fd_sc_hd__buf_8 repeater513 (.A(net56),
    .X(net513));
 sky130_fd_sc_hd__buf_8 repeater514 (.A(net45),
    .X(net514));
 sky130_fd_sc_hd__buf_8 repeater515 (.A(net43),
    .X(net515));
 sky130_fd_sc_hd__buf_8 repeater516 (.A(net39),
    .X(net516));
 sky130_fd_sc_hd__buf_8 repeater517 (.A(net36),
    .X(net517));
 sky130_fd_sc_hd__buf_8 repeater518 (.A(net30),
    .X(net518));
 sky130_fd_sc_hd__buf_8 repeater519 (.A(net25),
    .X(net519));
 sky130_fd_sc_hd__buf_8 repeater520 (.A(net21),
    .X(net520));
 sky130_fd_sc_hd__buf_8 repeater521 (.A(net20),
    .X(net521));
 sky130_fd_sc_hd__buf_8 repeater522 (.A(net2),
    .X(net522));
 sky130_fd_sc_hd__buf_8 repeater523 (.A(net14),
    .X(net523));
 sky130_fd_sc_hd__buf_8 repeater524 (.A(net13),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_17_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_21_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_20_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_22_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_26_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_23_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_opt_7_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_opt_8_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_opt_13_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_opt_9_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_29_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_opt_10_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_28_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_27_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_24_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_25_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_opt_12_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_opt_14_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_31_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_30_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_opt_1_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_opt_2_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_opt_4_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_opt_5_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_opt_6_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_7_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_13_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_15_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_14_0_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_5_10_0_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_11_0_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_8_0_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_9_0_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_opt_0_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_12_0_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_6_0_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_5_0_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_4_0_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_3_0_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_2_0_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_0_0_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_1_0_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_19_0_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_253_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk (.A(clknet_5_18_0_clk),
    .X(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk (.A(clknet_5_16_0_clk),
    .X(clknet_leaf_267_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_0_0_clk (.A(clknet_0_clk),
    .X(clknet_1_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_0_1_clk (.A(clknet_1_0_0_clk),
    .X(clknet_1_0_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_1_0_clk (.A(clknet_0_clk),
    .X(clknet_1_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_1_1_1_clk (.A(clknet_1_1_0_clk),
    .X(clknet_1_1_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_0_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_0_1_clk (.A(clknet_2_0_0_clk),
    .X(clknet_2_0_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_1_0_clk (.A(clknet_1_0_1_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_1_1_clk (.A(clknet_2_1_0_clk),
    .X(clknet_2_1_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_2_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_2_1_clk (.A(clknet_2_2_0_clk),
    .X(clknet_2_2_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_3_0_clk (.A(clknet_1_1_1_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_2_3_1_clk (.A(clknet_2_3_0_clk),
    .X(clknet_2_3_1_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_0_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_1_0_clk (.A(clknet_2_0_1_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_2_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_3_0_clk (.A(clknet_2_1_1_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_4_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_5_0_clk (.A(clknet_2_2_1_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_6_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_3_7_0_clk (.A(clknet_2_3_1_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_0_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_1_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_2_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_3_0_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_4_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_5_0_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_6_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_7_0_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_8_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_9_0_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_10_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_11_0_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_12_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_13_0_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_14_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_4_15_0_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_0_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_1_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_2_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_3_0_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_4_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_5_0_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_6_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_7_0_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_8_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_9_0_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_10_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_11_0_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_12_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_13_0_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_14_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_15_0_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_16_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_17_0_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_18_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_19_0_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_20_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_21_0_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_22_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_23_0_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_24_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_25_0_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_26_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_27_0_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_28_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_29_0_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_30_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30_0_clk));
 sky130_fd_sc_hd__clkbuf_2 clkbuf_5_31_0_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_0_clk (.A(clknet_5_5_0_clk),
    .X(clknet_opt_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_clk (.A(clknet_5_7_0_clk),
    .X(clknet_opt_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_clk (.A(clknet_5_7_0_clk),
    .X(clknet_opt_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_clk (.A(clknet_5_7_0_clk),
    .X(clknet_opt_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_clk (.A(clknet_5_7_0_clk),
    .X(clknet_opt_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_5_clk (.A(clknet_5_13_0_clk),
    .X(clknet_opt_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_6_clk (.A(clknet_5_15_0_clk),
    .X(clknet_opt_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_7_clk (.A(clknet_5_26_0_clk),
    .X(clknet_opt_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_8_clk (.A(clknet_5_27_0_clk),
    .X(clknet_opt_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_9_clk (.A(clknet_5_28_0_clk),
    .X(clknet_opt_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_10_clk (.A(clknet_5_29_0_clk),
    .X(clknet_opt_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_11_clk (.A(clknet_5_29_0_clk),
    .X(clknet_opt_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_12_clk (.A(clknet_5_29_0_clk),
    .X(clknet_opt_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_13_clk (.A(clknet_5_30_0_clk),
    .X(clknet_opt_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_14_clk (.A(clknet_5_31_0_clk),
    .X(clknet_opt_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_15_clk (.A(clknet_5_31_0_clk),
    .X(clknet_opt_15_clk));
endmodule
